// Benchmark "c7552" written by ABC on Wed Oct 05 14:38:34 2022

module c7552 ( 
    \1 , 5, 9, 12, 15, 18, 23, 26, 29, 32, 35, 38, 41, 44, 47, 50, 53, 54,
    55, 56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 69, 70, 73, 74, 75, 76,
    77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 94, 97, 100, 103,
    106, 109, 110, 111, 112, 113, 114, 115, 118, 121, 124, 127, 130, 133,
    134, 135, 138, 141, 144, 147, 150, 151, 152, 153, 154, 155, 156, 157,
    158, 159, 160, 161, 162, 163, 164, 165, 166, 167, 168, 169, 170, 171,
    172, 173, 174, 175, 176, 177, 178, 179, 180, 181, 182, 183, 184, 185,
    186, 187, 188, 189, 190, 191, 192, 193, 194, 195, 196, 197, 198, 199,
    200, 201, 202, 203, 204, 205, 206, 207, 208, 209, 210, 211, 212, 213,
    214, 215, 216, 217, 218, 219, 220, 221, 222, 223, 224, 225, 226, 227,
    228, 229, 230, 231, 232, 233, 234, 235, 236, 237, 238, 239, 240, 241,
    242, 245, 248, 251, 254, 257, 260, 263, 267, 271, 274, 277, 280, 283,
    286, 289, 293, 296, 299, 303, 307, 310, 313, 316, 319, 322, 325, 328,
    331, 334, 337, 340, 343, 346, 349, 352, 355, 358, 361, 364, 367, 382,
    387, 388, 478, 482, 484, 486, 489, 492, 501, 505, 507, 509, 511, 513,
    515, 517, 519, 535, 537, 539, 541, 543, 545, 547, 549, 551, 553, 556,
    559, 561, 563, 565, 567, 569, 571, 573, 582, 643, 707, 813, 881, 882,
    883, 884, 885, 889, 945, 1110, 1111, 1112, 1113, 1114, 1489, 1490,
    1781, 10025, 10101, 10102, 10103, 10104, 10109, 10110, 10111, 10112,
    10350, 10351, 10352, 10353, 10574, 10575, 10576, 10628, 10632, 10641,
    10704, 10706, 10711, 10712, 10713, 10714, 10715, 10716, 10717, 10718,
    10729, 10759, 10760, 10761, 10762, 10763, 10827, 10837, 10838, 10839,
    10840, 10868, 10869, 10870, 10871, 10905, 10906, 10907, 10908, 11333,
    11334, 11340, 11342  );
  input  \1 , 5, 9, 12, 15, 18, 23, 26, 29, 32, 35, 38, 41, 44, 47, 50,
    53, 54, 55, 56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 69, 70, 73, 74,
    75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 94, 97,
    100, 103, 106, 109, 110, 111, 112, 113, 114, 115, 118, 121, 124, 127,
    130, 133, 134, 135, 138, 141, 144, 147, 150, 151, 152, 153, 154, 155,
    156, 157, 158, 159, 160, 161, 162, 163, 164, 165, 166, 167, 168, 169,
    170, 171, 172, 173, 174, 175, 176, 177, 178, 179, 180, 181, 182, 183,
    184, 185, 186, 187, 188, 189, 190, 191, 192, 193, 194, 195, 196, 197,
    198, 199, 200, 201, 202, 203, 204, 205, 206, 207, 208, 209, 210, 211,
    212, 213, 214, 215, 216, 217, 218, 219, 220, 221, 222, 223, 224, 225,
    226, 227, 228, 229, 230, 231, 232, 233, 234, 235, 236, 237, 238, 239,
    240, 241, 242, 245, 248, 251, 254, 257, 260, 263, 267, 271, 274, 277,
    280, 283, 286, 289, 293, 296, 299, 303, 307, 310, 313, 316, 319, 322,
    325, 328, 331, 334, 337, 340, 343, 346, 349, 352, 355, 358, 361, 364,
    367, 382;
  output 387, 388, 478, 482, 484, 486, 489, 492, 501, 505, 507, 509, 511, 513,
    515, 517, 519, 535, 537, 539, 541, 543, 545, 547, 549, 551, 553, 556,
    559, 561, 563, 565, 567, 569, 571, 573, 582, 643, 707, 813, 881, 882,
    883, 884, 885, 889, 945, 1110, 1111, 1112, 1113, 1114, 1489, 1490,
    1781, 10025, 10101, 10102, 10103, 10104, 10109, 10110, 10111, 10112,
    10350, 10351, 10352, 10353, 10574, 10575, 10576, 10628, 10632, 10641,
    10704, 10706, 10711, 10712, 10713, 10714, 10715, 10716, 10717, 10718,
    10729, 10759, 10760, 10761, 10762, 10763, 10827, 10837, 10838, 10839,
    10840, 10868, 10869, 10870, 10871, 10905, 10906, 10907, 10908, 11333,
    11334, 11340, 11342;
  wire n321, n325, n326, n327, n328, n329, n331, n332, n333, n334, n335,
    n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
    n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
    n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
    n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
    n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
    n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
    n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
    n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
    n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
    n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
    n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
    n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
    n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
    n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
    n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
    n516, n517, n518, n519, n520, n521, n522, n523, n525, n526, n527, n528,
    n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
    n541, n542, n543, n544, n545, n546, n547, n548, n549, n551, n552, n553,
    n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
    n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
    n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
    n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
    n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
    n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
    n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
    n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
    n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
    n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
    n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
    n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
    n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
    n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
    n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
    n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
    n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
    n758, n759, n760, n761, n762, n763, n764, n768, n774, n787, n788, n789,
    n790, n791, n792, n794, n795, n796, n797, n798, n800, n801, n802, n804,
    n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n817, n818,
    n819, n820, n821, n822, n823, n825, n826, n827, n830, n831, n832, n833,
    n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
    n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
    n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
    n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
    n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n893, n894,
    n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
    n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
    n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
    n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
    n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
    n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n967,
    n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
    n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
    n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
    n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
    n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
    n1023, n1024, n1025, n1026, n1027, n1028, n1030, n1031, n1032, n1034,
    n1035, n1036, n1038, n1039, n1041, n1042, n1043, n1044, n1045, n1046,
    n1048, n1049, n1050, n1053, n1055, n1056, n1057, n1058, n1059, n1060,
    n1061, n1063, n1064, n1065, n1066, n1068, n1069, n1070, n1071, n1073,
    n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1083, n1084, n1085,
    n1086, n1087, n1089, n1090, n1091, n1092, n1094, n1096, n1101, n1102,
    n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
    n1114, n1115, n1116, n1117, n1119, n1120, n1121, n1123, n1125, n1126,
    n1128, n1129, n1130, n1131, n1134, n1135, n1136, n1137, n1138, n1139,
    n1140, n1142, n1143, n1144, n1145, n1147, n1148, n1149, n1150, n1152,
    n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1164, n1165,
    n1166, n1167, n1168, n1170, n1171, n1172, n1175, n1176, n1177, n1178,
    n1179, n1180, n1181, n1182, n1185, n1187, n1188, n1189, n1190, n1191,
    n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
    n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
    n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1221, n1222,
    n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
    n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
    n1243, n1244, n1245, n1248, n1249, n1250, n1251, n1252, n1253, n1255,
    n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
    n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
    n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
    n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
    n1296, n1297, n1298, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
    n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
    n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
    n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
    n1337, n1338, n1339, n1340, n1341, n1342;
  INV_X1    g0000(.A(15), .ZN(582));
  OR2_X1    g0001(.A1(57), .A2(5), .ZN(881));
  NAND4_X1  g0002(.A1(228), .A2(184), .A3(150), .A4(240), .ZN(882));
  NAND4_X1  g0003(.A1(218), .A2(210), .A3(152), .A4(230), .ZN(883));
  NAND4_X1  g0004(.A1(185), .A2(183), .A3(182), .A4(186), .ZN(884));
  NAND4_X1  g0005(.A1(188), .A2(172), .A3(162), .A4(199), .ZN(885));
  INV_X1    g0006(.A(5), .ZN(n321));
  NAND2_X1  g0007(.A1(242), .A2(n321), .ZN(1110));
  NAND3_X1  g0008(.A1(134), .A2(133), .A3(n321), .ZN(1113));
  AND2_X1   g0009(.A1(163), .A2(\1 ), .ZN(1781));
  INV_X1    g0010(.A(18), .ZN(n325));
  NAND2_X1  g0011(.A1(41), .A2(n325), .ZN(n326));
  INV_X1    g0012(.A(310), .ZN(n327));
  NOR2_X1   g0013(.A1(n327), .A2(18), .ZN(n328));
  XNOR2_X1  g0014(.A(n328), .B(n326), .ZN(n329));
  XNOR2_X1  g0015(.A(n329), .B(367), .ZN(10025));
  INV_X1    g0016(.A(38), .ZN(n331));
  AND2_X1   g0017(.A1(382), .A2(267), .ZN(n332));
  XNOR2_X1  g0018(.A(n332), .B(n331), .ZN(n333));
  AND2_X1   g0019(.A1(382), .A2(263), .ZN(n334));
  XNOR2_X1  g0020(.A(n334), .B(n331), .ZN(n335));
  NOR2_X1   g0021(.A1(n335), .A2(n333), .ZN(n336));
  INV_X1    g0022(.A(254), .ZN(n337));
  INV_X1    g0023(.A(216), .ZN(n338));
  AOI22_X1  g0024(.A1(18), .A2(n338), .B1(12), .B2(9), .ZN(n339));
  XNOR2_X1  g0025(.A(n339), .B(n337), .ZN(n340));
  INV_X1    g0026(.A(251), .ZN(n341));
  INV_X1    g0027(.A(209), .ZN(n342));
  AOI22_X1  g0028(.A1(18), .A2(n342), .B1(12), .B2(9), .ZN(n343));
  XNOR2_X1  g0029(.A(n343), .B(n341), .ZN(n344));
  NOR2_X1   g0030(.A1(n344), .A2(n340), .ZN(n345));
  NAND2_X1  g0031(.A1(12), .A2(9), .ZN(n346));
  OAI21_X1  g0032(.A(n346), .B1(213), .B2(n325), .ZN(n347));
  XNOR2_X1  g0033(.A(n347), .B(260), .ZN(n348));
  INV_X1    g0034(.A(n348), .ZN(n349));
  INV_X1    g0035(.A(215), .ZN(n350));
  AOI22_X1  g0036(.A1(18), .A2(n350), .B1(12), .B2(9), .ZN(n351));
  XNOR2_X1  g0037(.A(n351), .B(106), .ZN(n352));
  INV_X1    g0038(.A(214), .ZN(n353));
  AOI22_X1  g0039(.A1(18), .A2(n353), .B1(12), .B2(9), .ZN(n354));
  XNOR2_X1  g0040(.A(n354), .B(257), .ZN(n355));
  AND4_X1   g0041(.A1(n352), .A2(n349), .A3(n345), .A4(n355), .ZN(n356));
  AND2_X1   g0042(.A1(n356), .A2(n336), .ZN(n357));
  INV_X1    g0043(.A(303), .ZN(n358));
  INV_X1    g0044(.A(153), .ZN(n359));
  AOI22_X1  g0045(.A1(18), .A2(n359), .B1(12), .B2(9), .ZN(n360));
  XNOR2_X1  g0046(.A(n360), .B(n358), .ZN(n361));
  INV_X1    g0047(.A(n361), .ZN(n362));
  INV_X1    g0048(.A(156), .ZN(n363));
  AOI22_X1  g0049(.A1(18), .A2(n363), .B1(12), .B2(9), .ZN(n364));
  XNOR2_X1  g0050(.A(n364), .B(293), .ZN(n365));
  INV_X1    g0051(.A(155), .ZN(n366));
  AOI22_X1  g0052(.A1(18), .A2(n366), .B1(12), .B2(9), .ZN(n367));
  XNOR2_X1  g0053(.A(n367), .B(296), .ZN(n368));
  INV_X1    g0054(.A(299), .ZN(n369));
  INV_X1    g0055(.A(154), .ZN(n370));
  AOI22_X1  g0056(.A1(18), .A2(n370), .B1(12), .B2(9), .ZN(n371));
  XNOR2_X1  g0057(.A(n371), .B(n369), .ZN(n372));
  INV_X1    g0058(.A(n372), .ZN(n373));
  NAND4_X1  g0059(.A1(n368), .A2(n365), .A3(n362), .A4(n373), .ZN(n374));
  INV_X1    g0060(.A(289), .ZN(n375));
  INV_X1    g0061(.A(157), .ZN(n376));
  AOI22_X1  g0062(.A1(18), .A2(n376), .B1(12), .B2(9), .ZN(n377));
  XNOR2_X1  g0063(.A(n377), .B(n375), .ZN(n378));
  INV_X1    g0064(.A(n378), .ZN(n379));
  INV_X1    g0065(.A(280), .ZN(n380));
  MUX2_X1   g0066(.S(18), .B(160), .A(138), .ZN(n381));
  XNOR2_X1  g0067(.A(n381), .B(n380), .ZN(n382));
  INV_X1    g0068(.A(277), .ZN(n383));
  MUX2_X1   g0069(.S(18), .B(151), .A(147), .ZN(n384));
  XNOR2_X1  g0070(.A(n384), .B(n383), .ZN(n385));
  NOR2_X1   g0071(.A1(n385), .A2(n382), .ZN(n386));
  INV_X1    g0072(.A(283), .ZN(n387));
  MUX2_X1   g0073(.S(18), .B(159), .A(144), .ZN(n388));
  XNOR2_X1  g0074(.A(n388), .B(n387), .ZN(n389));
  INV_X1    g0075(.A(n389), .ZN(n390));
  INV_X1    g0076(.A(286), .ZN(n391));
  MUX2_X1   g0077(.S(18), .B(158), .A(135), .ZN(n392));
  XNOR2_X1  g0078(.A(n392), .B(n391), .ZN(n393));
  INV_X1    g0079(.A(n393), .ZN(n394));
  NAND4_X1  g0080(.A1(n390), .A2(n386), .A3(n379), .A4(n394), .ZN(n395));
  NOR2_X1   g0081(.A1(n395), .A2(n374), .ZN(n396));
  INV_X1    g0082(.A(364), .ZN(n397));
  MUX2_X1   g0083(.S(18), .B(219), .A(66), .ZN(n398));
  XNOR2_X1  g0084(.A(n398), .B(n397), .ZN(n399));
  INV_X1    g0085(.A(355), .ZN(n400));
  MUX2_X1   g0086(.S(18), .B(222), .A(35), .ZN(n401));
  XNOR2_X1  g0087(.A(n401), .B(n400), .ZN(n402));
  INV_X1    g0088(.A(358), .ZN(n403));
  MUX2_X1   g0089(.S(18), .B(221), .A(32), .ZN(n404));
  XNOR2_X1  g0090(.A(n404), .B(n403), .ZN(n405));
  INV_X1    g0091(.A(361), .ZN(n406));
  MUX2_X1   g0092(.S(18), .B(220), .A(50), .ZN(n407));
  XNOR2_X1  g0093(.A(n407), .B(n406), .ZN(n408));
  NOR4_X1   g0094(.A1(n405), .A2(n402), .A3(n399), .A4(n408), .ZN(n409));
  INV_X1    g0095(.A(343), .ZN(n410));
  MUX2_X1   g0096(.S(18), .B(226), .A(97), .ZN(n411));
  XNOR2_X1  g0097(.A(n411), .B(n410), .ZN(n412));
  INV_X1    g0098(.A(340), .ZN(n413));
  MUX2_X1   g0099(.S(18), .B(217), .A(118), .ZN(n414));
  XNOR2_X1  g0100(.A(n414), .B(n413), .ZN(n415));
  OR2_X1    g0101(.A1(n415), .A2(n412), .ZN(n416));
  INV_X1    g0102(.A(352), .ZN(n417));
  MUX2_X1   g0103(.S(18), .B(223), .A(47), .ZN(n418));
  XNOR2_X1  g0104(.A(n418), .B(n417), .ZN(n419));
  INV_X1    g0105(.A(346), .ZN(n420));
  MUX2_X1   g0106(.S(18), .B(225), .A(94), .ZN(n421));
  XNOR2_X1  g0107(.A(n421), .B(n420), .ZN(n422));
  INV_X1    g0108(.A(349), .ZN(n423));
  MUX2_X1   g0109(.S(18), .B(224), .A(121), .ZN(n424));
  XNOR2_X1  g0110(.A(n424), .B(n423), .ZN(n425));
  NOR4_X1   g0111(.A1(n422), .A2(n419), .A3(n416), .A4(n425), .ZN(n426));
  AND2_X1   g0112(.A1(n426), .A2(n409), .ZN(n427));
  INV_X1    g0113(.A(334), .ZN(n428));
  MUX2_X1   g0114(.S(18), .B(231), .A(100), .ZN(n429));
  XNOR2_X1  g0115(.A(n429), .B(n428), .ZN(n430));
  INV_X1    g0116(.A(331), .ZN(n431));
  MUX2_X1   g0117(.S(18), .B(232), .A(124), .ZN(n432));
  XNOR2_X1  g0118(.A(n432), .B(n431), .ZN(n433));
  INV_X1    g0119(.A(328), .ZN(n434));
  MUX2_X1   g0120(.S(18), .B(233), .A(127), .ZN(n435));
  AND2_X1   g0121(.A1(n435), .A2(n434), .ZN(n436));
  INV_X1    g0122(.A(n436), .ZN(n437));
  NOR3_X1   g0123(.A1(n437), .A2(n433), .A3(n430), .ZN(n438));
  INV_X1    g0124(.A(325), .ZN(n439));
  MUX2_X1   g0125(.S(18), .B(234), .A(130), .ZN(n440));
  AND2_X1   g0126(.A1(n440), .A2(n439), .ZN(n441));
  INV_X1    g0127(.A(n441), .ZN(n442));
  XNOR2_X1  g0128(.A(n435), .B(n434), .ZN(n443));
  NOR4_X1   g0129(.A1(n442), .A2(n433), .A3(n430), .A4(n443), .ZN(n444));
  NAND2_X1  g0130(.A1(n429), .A2(n428), .ZN(n445));
  NAND2_X1  g0131(.A1(n432), .A2(n431), .ZN(n446));
  OAI21_X1  g0132(.A(n445), .B1(n446), .B2(n430), .ZN(n447));
  NOR3_X1   g0133(.A1(n447), .A2(n444), .A3(n438), .ZN(n448));
  XNOR2_X1  g0134(.A(n440), .B(n439), .ZN(n449));
  OR4_X1    g0135(.A1(n443), .A2(n433), .A3(n430), .A4(n449), .ZN(n450));
  INV_X1    g0136(.A(313), .ZN(n451));
  MUX2_X1   g0137(.S(18), .B(238), .A(29), .ZN(n452));
  XNOR2_X1  g0138(.A(n452), .B(n451), .ZN(n453));
  INV_X1    g0139(.A(316), .ZN(n454));
  MUX2_X1   g0140(.S(18), .B(237), .A(26), .ZN(n455));
  XNOR2_X1  g0141(.A(n455), .B(n454), .ZN(n456));
  OR2_X1    g0142(.A1(n456), .A2(n453), .ZN(n457));
  INV_X1    g0143(.A(322), .ZN(n458));
  MUX2_X1   g0144(.S(18), .B(235), .A(103), .ZN(n459));
  XNOR2_X1  g0145(.A(n459), .B(n458), .ZN(n460));
  INV_X1    g0146(.A(319), .ZN(n461));
  MUX2_X1   g0147(.S(18), .B(236), .A(23), .ZN(n462));
  XNOR2_X1  g0148(.A(n462), .B(n461), .ZN(n463));
  MUX2_X1   g0149(.S(18), .B(229), .A(41), .ZN(n464));
  NAND3_X1  g0150(.A1(n464), .A2(n327), .A3(n325), .ZN(n465));
  NOR4_X1   g0151(.A1(n463), .A2(n460), .A3(n457), .A4(n465), .ZN(n466));
  INV_X1    g0152(.A(n463), .ZN(n467));
  NAND3_X1  g0153(.A1(n467), .A2(n455), .A3(n454), .ZN(n468));
  NAND2_X1  g0154(.A1(n452), .A2(n451), .ZN(n469));
  NOR4_X1   g0155(.A1(n463), .A2(n460), .A3(n456), .A4(n469), .ZN(n470));
  NAND2_X1  g0156(.A1(n462), .A2(n461), .ZN(n471));
  NOR2_X1   g0157(.A1(n471), .A2(n460), .ZN(n472));
  AOI211_X1 g0158(.A(n470), .B(n472), .C1(n459), .C2(n458), .ZN(n473));
  OAI21_X1  g0159(.A(n473), .B1(n468), .B2(n460), .ZN(n474));
  NOR2_X1   g0160(.A1(n474), .A2(n466), .ZN(n475));
  OAI21_X1  g0161(.A(n448), .B1(n475), .B2(n450), .ZN(n476));
  NAND4_X1  g0162(.A1(n427), .A2(n396), .A3(n357), .A4(n476), .ZN(n477));
  AND2_X1   g0163(.A1(n404), .A2(n403), .ZN(n478));
  INV_X1    g0164(.A(n478), .ZN(n479));
  OR3_X1    g0165(.A1(n479), .A2(n408), .A3(n399), .ZN(n480));
  INV_X1    g0166(.A(n399), .ZN(n481));
  INV_X1    g0167(.A(n405), .ZN(n482));
  INV_X1    g0168(.A(n408), .ZN(n483));
  AND2_X1   g0169(.A1(n401), .A2(n400), .ZN(n484));
  NAND4_X1  g0170(.A1(n483), .A2(n482), .A3(n481), .A4(n484), .ZN(n485));
  AND2_X1   g0171(.A1(n398), .A2(n397), .ZN(n486));
  AND2_X1   g0172(.A1(n407), .A2(n406), .ZN(n487));
  AOI21_X1  g0173(.A(n486), .B1(n487), .B2(n481), .ZN(n488));
  NAND3_X1  g0174(.A1(n488), .A2(n485), .A3(n480), .ZN(n489));
  INV_X1    g0175(.A(n419), .ZN(n490));
  INV_X1    g0176(.A(n425), .ZN(n491));
  NOR2_X1   g0177(.A1(n422), .A2(n412), .ZN(n492));
  AND2_X1   g0178(.A1(n414), .A2(n413), .ZN(n493));
  NAND4_X1  g0179(.A1(n492), .A2(n491), .A3(n490), .A4(n493), .ZN(n494));
  NAND4_X1  g0180(.A1(n421), .A2(n490), .A3(n420), .A4(n491), .ZN(n495));
  NAND2_X1  g0181(.A1(n411), .A2(n410), .ZN(n496));
  OR4_X1    g0182(.A1(n425), .A2(n422), .A3(n419), .A4(n496), .ZN(n497));
  AND2_X1   g0183(.A1(n418), .A2(n417), .ZN(n498));
  AND2_X1   g0184(.A1(n424), .A2(n423), .ZN(n499));
  AOI21_X1  g0185(.A(n498), .B1(n499), .B2(n490), .ZN(n500));
  NAND4_X1  g0186(.A1(n497), .A2(n495), .A3(n494), .A4(n500), .ZN(n501));
  AOI21_X1  g0187(.A(n489), .B1(n501), .B2(n409), .ZN(n502));
  NOR3_X1   g0188(.A1(n502), .A2(n395), .A3(n374), .ZN(n503));
  NAND2_X1  g0189(.A1(n503), .A2(n357), .ZN(n504));
  AOI21_X1  g0190(.A(n331), .B1(n334), .B2(n332), .ZN(n505));
  INV_X1    g0191(.A(106), .ZN(n506));
  XNOR2_X1  g0192(.A(n351), .B(n506), .ZN(n507));
  NOR2_X1   g0193(.A1(n507), .A2(n340), .ZN(n508));
  AOI221_X1 g0194(.A(251), .B1(18), .B2(n342), .C1(12), .C2(9), .ZN(n509));
  AND4_X1   g0195(.A1(n508), .A2(n355), .A3(n349), .A4(n509), .ZN(n510));
  INV_X1    g0196(.A(257), .ZN(n511));
  XNOR2_X1  g0197(.A(n354), .B(n511), .ZN(n512));
  OAI211_X1 g0198(.A(n506), .B(n346), .C1(215), .C2(n325), .ZN(n513));
  NOR3_X1   g0199(.A1(n513), .A2(n512), .A3(n348), .ZN(n514));
  OAI211_X1 g0200(.A(n337), .B(n346), .C1(216), .C2(n325), .ZN(n515));
  NOR4_X1   g0201(.A1(n512), .A2(n507), .A3(n348), .A4(n515), .ZN(n516));
  NOR2_X1   g0202(.A1(n347), .A2(260), .ZN(n517));
  AOI221_X1 g0203(.A(257), .B1(18), .B2(n353), .C1(12), .C2(9), .ZN(n518));
  AOI211_X1 g0204(.A(n517), .B(n516), .C1(n349), .C2(n518), .ZN(n519));
  INV_X1    g0205(.A(n519), .ZN(n520));
  NOR3_X1   g0206(.A1(n520), .A2(n514), .A3(n510), .ZN(n521));
  INV_X1    g0207(.A(n521), .ZN(n522));
  AOI21_X1  g0208(.A(n505), .B1(n522), .B2(n336), .ZN(n523));
  OR2_X1    g0209(.A1(n460), .A2(n456), .ZN(n525));
  NOR4_X1   g0210(.A1(n463), .A2(n453), .A3(n329), .A4(n525), .ZN(n526));
  NAND4_X1  g0211(.A1(n774), .A2(n427), .A3(367), .A4(n526), .ZN(n527));
  NOR3_X1   g0212(.A1(n527), .A2(n395), .A3(n374), .ZN(n528));
  AOI221_X1 g0213(.A(296), .B1(18), .B2(n366), .C1(12), .C2(9), .ZN(n529));
  NAND3_X1  g0214(.A1(n529), .A2(n373), .A3(n362), .ZN(n530));
  AOI221_X1 g0215(.A(293), .B1(18), .B2(n363), .C1(12), .C2(9), .ZN(n531));
  NAND4_X1  g0216(.A1(n373), .A2(n368), .A3(n362), .A4(n531), .ZN(n532));
  AOI221_X1 g0217(.A(303), .B1(18), .B2(n359), .C1(12), .C2(9), .ZN(n533));
  AOI221_X1 g0218(.A(299), .B1(18), .B2(n370), .C1(12), .C2(9), .ZN(n534));
  AOI21_X1  g0219(.A(n533), .B1(n534), .B2(n362), .ZN(n535));
  AND3_X1   g0220(.A1(n535), .A2(n532), .A3(n530), .ZN(n536));
  AND2_X1   g0221(.A1(n392), .A2(n391), .ZN(n537));
  AND2_X1   g0222(.A1(n537), .A2(n379), .ZN(n538));
  NAND3_X1  g0223(.A1(n394), .A2(n388), .A3(n387), .ZN(n539));
  OAI211_X1 g0224(.A(n375), .B(n346), .C1(157), .C2(n325), .ZN(n540));
  OAI21_X1  g0225(.A(n540), .B1(n539), .B2(n378), .ZN(n541));
  NOR2_X1   g0226(.A1(n389), .A2(n382), .ZN(n542));
  AND2_X1   g0227(.A1(n384), .A2(n383), .ZN(n543));
  AND4_X1   g0228(.A1(n542), .A2(n394), .A3(n379), .A4(n543), .ZN(n544));
  NAND2_X1  g0229(.A1(n381), .A2(n380), .ZN(n545));
  NOR4_X1   g0230(.A1(n393), .A2(n389), .A3(n378), .A4(n545), .ZN(n546));
  NOR4_X1   g0231(.A1(n544), .A2(n541), .A3(n538), .A4(n546), .ZN(n547));
  OAI21_X1  g0232(.A(n536), .B1(n547), .B2(n374), .ZN(n548));
  OAI21_X1  g0233(.A(n357), .B1(n548), .B2(n528), .ZN(n549));
  NAND4_X1  g0234(.A1(n523), .A2(n504), .A3(n477), .A4(n549), .ZN(10101));
  INV_X1    g0235(.A(382), .ZN(n551));
  NOR2_X1   g0236(.A1(n551), .A2(271), .ZN(n552));
  XNOR2_X1  g0237(.A(n552), .B(n331), .ZN(n553));
  NOR2_X1   g0238(.A1(n551), .A2(245), .ZN(n554));
  XNOR2_X1  g0239(.A(n554), .B(n331), .ZN(n555));
  INV_X1    g0240(.A(88), .ZN(n556));
  MUX2_X1   g0241(.S(18), .B(260), .A(n556), .ZN(n557));
  OAI21_X1  g0242(.A(n346), .B1(166), .B2(n325), .ZN(n558));
  XNOR2_X1  g0243(.A(n558), .B(n557), .ZN(n559));
  INV_X1    g0244(.A(n559), .ZN(n560));
  MUX2_X1   g0245(.S(18), .B(n341), .A(113), .ZN(n561));
  XOR2_X1   g0246(.A(n561), .B(n346), .ZN(n562));
  MUX2_X1   g0247(.S(18), .B(n511), .A(112), .ZN(n563));
  OAI21_X1  g0248(.A(n346), .B1(167), .B2(n325), .ZN(n564));
  XOR2_X1   g0249(.A(n564), .B(n563), .ZN(n565));
  MUX2_X1   g0250(.S(18), .B(n506), .A(87), .ZN(n566));
  OAI21_X1  g0251(.A(n346), .B1(168), .B2(n325), .ZN(n567));
  XOR2_X1   g0252(.A(n567), .B(n566), .ZN(n568));
  MUX2_X1   g0253(.S(18), .B(n337), .A(111), .ZN(n569));
  OAI21_X1  g0254(.A(n346), .B1(169), .B2(n325), .ZN(n570));
  XOR2_X1   g0255(.A(n570), .B(n569), .ZN(n571));
  NOR3_X1   g0256(.A1(n571), .A2(n568), .A3(n565), .ZN(n572));
  NAND3_X1  g0257(.A1(n572), .A2(n562), .A3(n560), .ZN(n573));
  NOR3_X1   g0258(.A1(n573), .A2(n555), .A3(n553), .ZN(n574));
  MUX2_X1   g0259(.S(18), .B(n358), .A(110), .ZN(n575));
  INV_X1    g0260(.A(173), .ZN(n576));
  AOI22_X1  g0261(.A1(18), .A2(n576), .B1(12), .B2(9), .ZN(n577));
  XNOR2_X1  g0262(.A(n577), .B(n575), .ZN(n578));
  INV_X1    g0263(.A(293), .ZN(n579));
  MUX2_X1   g0264(.S(18), .B(n579), .A(63), .ZN(n580));
  OAI21_X1  g0265(.A(n346), .B1(176), .B2(n325), .ZN(n581));
  XOR2_X1   g0266(.A(n581), .B(n580), .ZN(n582));
  MUX2_X1   g0267(.S(18), .B(n369), .A(109), .ZN(n583));
  OAI21_X1  g0268(.A(n346), .B1(174), .B2(n325), .ZN(n584));
  XOR2_X1   g0269(.A(n584), .B(n583), .ZN(n585));
  INV_X1    g0270(.A(296), .ZN(n586));
  MUX2_X1   g0271(.S(18), .B(n586), .A(86), .ZN(n587));
  INV_X1    g0272(.A(175), .ZN(n588));
  AOI22_X1  g0273(.A1(18), .A2(n588), .B1(12), .B2(9), .ZN(n589));
  XNOR2_X1  g0274(.A(n589), .B(n587), .ZN(n590));
  OR4_X1    g0275(.A1(n585), .A2(n582), .A3(n578), .A4(n590), .ZN(n591));
  MUX2_X1   g0276(.S(18), .B(n375), .A(64), .ZN(n592));
  OAI21_X1  g0277(.A(n346), .B1(177), .B2(n325), .ZN(n593));
  XOR2_X1   g0278(.A(n593), .B(n592), .ZN(n594));
  MUX2_X1   g0279(.S(18), .B(n391), .A(85), .ZN(n595));
  INV_X1    g0280(.A(n595), .ZN(n596));
  AND2_X1   g0281(.A1(178), .A2(18), .ZN(n597));
  AOI21_X1  g0282(.A(n597), .B1(135), .B2(n325), .ZN(n598));
  NOR3_X1   g0283(.A1(n598), .A2(n596), .A3(n594), .ZN(n599));
  XOR2_X1   g0284(.A(n598), .B(n595), .ZN(n600));
  INV_X1    g0285(.A(84), .ZN(n601));
  MUX2_X1   g0286(.S(18), .B(283), .A(n601), .ZN(n602));
  MUX2_X1   g0287(.S(18), .B(179), .A(144), .ZN(n603));
  INV_X1    g0288(.A(n603), .ZN(n604));
  NOR4_X1   g0289(.A1(n602), .A2(n600), .A3(n594), .A4(n604), .ZN(n605));
  OR2_X1    g0290(.A1(177), .A2(n325), .ZN(n606));
  AND3_X1   g0291(.A1(n606), .A2(n592), .A3(n346), .ZN(n607));
  XNOR2_X1  g0292(.A(n604), .B(n602), .ZN(n608));
  INV_X1    g0293(.A(83), .ZN(n609));
  MUX2_X1   g0294(.S(18), .B(280), .A(n609), .ZN(n610));
  MUX2_X1   g0295(.S(18), .B(180), .A(138), .ZN(n611));
  INV_X1    g0296(.A(n611), .ZN(n612));
  XNOR2_X1  g0297(.A(n612), .B(n610), .ZN(n613));
  MUX2_X1   g0298(.S(18), .B(n383), .A(65), .ZN(n614));
  MUX2_X1   g0299(.S(18), .B(171), .A(147), .ZN(n615));
  NAND2_X1  g0300(.A1(n615), .A2(n614), .ZN(n616));
  OR4_X1    g0301(.A1(n613), .A2(n608), .A3(n600), .A4(n616), .ZN(n617));
  OR4_X1    g0302(.A1(n610), .A2(n608), .A3(n600), .A4(n612), .ZN(n618));
  AOI21_X1  g0303(.A(n594), .B1(n618), .B2(n617), .ZN(n619));
  NOR4_X1   g0304(.A1(n607), .A2(n605), .A3(n599), .A4(n619), .ZN(n620));
  NAND2_X1  g0305(.A1(n589), .A2(n587), .ZN(n621));
  OR3_X1    g0306(.A1(n621), .A2(n585), .A3(n578), .ZN(n622));
  OAI211_X1 g0307(.A(n346), .B(n580), .C1(176), .C2(n325), .ZN(n623));
  NOR4_X1   g0308(.A1(n590), .A2(n585), .A3(n578), .A4(n623), .ZN(n624));
  OAI211_X1 g0309(.A(n346), .B(n583), .C1(174), .C2(n325), .ZN(n625));
  NOR2_X1   g0310(.A1(n625), .A2(n578), .ZN(n626));
  AOI211_X1 g0311(.A(n624), .B(n626), .C1(n577), .C2(n575), .ZN(n627));
  OAI211_X1 g0312(.A(n622), .B(n627), .C1(n620), .C2(n591), .ZN(n628));
  NAND2_X1  g0313(.A1(n628), .A2(n574), .ZN(n629));
  NAND2_X1  g0314(.A1(n561), .A2(n346), .ZN(n630));
  OR3_X1    g0315(.A1(n571), .A2(n568), .A3(n559), .ZN(n631));
  NOR3_X1   g0316(.A1(n631), .A2(n630), .A3(n565), .ZN(n632));
  OAI211_X1 g0317(.A(n346), .B(n566), .C1(168), .C2(n325), .ZN(n633));
  NOR3_X1   g0318(.A1(n633), .A2(n565), .A3(n559), .ZN(n634));
  OAI211_X1 g0319(.A(n346), .B(n569), .C1(169), .C2(n325), .ZN(n635));
  NOR4_X1   g0320(.A1(n568), .A2(n565), .A3(n559), .A4(n635), .ZN(n636));
  OR2_X1    g0321(.A1(n558), .A2(n557), .ZN(n637));
  OAI211_X1 g0322(.A(n346), .B(n563), .C1(167), .C2(n325), .ZN(n638));
  OAI21_X1  g0323(.A(n637), .B1(n638), .B2(n559), .ZN(n639));
  NOR4_X1   g0324(.A1(n636), .A2(n634), .A3(n632), .A4(n639), .ZN(n640));
  NOR3_X1   g0325(.A1(n640), .A2(n555), .A3(n553), .ZN(n641));
  MUX2_X1   g0326(.S(18), .B(n397), .A(62), .ZN(n642));
  MUX2_X1   g0327(.S(18), .B(189), .A(66), .ZN(n643));
  XNOR2_X1  g0328(.A(n643), .B(n642), .ZN(n644));
  MUX2_X1   g0329(.S(18), .B(n400), .A(79), .ZN(n645));
  MUX2_X1   g0330(.S(18), .B(192), .A(35), .ZN(n646));
  XNOR2_X1  g0331(.A(n646), .B(n645), .ZN(n647));
  MUX2_X1   g0332(.S(18), .B(n406), .A(61), .ZN(n648));
  MUX2_X1   g0333(.S(18), .B(190), .A(50), .ZN(n649));
  XNOR2_X1  g0334(.A(n649), .B(n648), .ZN(n650));
  MUX2_X1   g0335(.S(18), .B(n403), .A(60), .ZN(n651));
  MUX2_X1   g0336(.S(18), .B(191), .A(32), .ZN(n652));
  XNOR2_X1  g0337(.A(n652), .B(n651), .ZN(n653));
  NOR4_X1   g0338(.A1(n650), .A2(n647), .A3(n644), .A4(n653), .ZN(n654));
  INV_X1    g0339(.A(80), .ZN(n655));
  MUX2_X1   g0340(.S(18), .B(352), .A(n655), .ZN(n656));
  MUX2_X1   g0341(.S(18), .B(193), .A(47), .ZN(n657));
  XOR2_X1   g0342(.A(n657), .B(n656), .ZN(n658));
  MUX2_X1   g0343(.S(18), .B(n413), .A(77), .ZN(n659));
  MUX2_X1   g0344(.S(18), .B(187), .A(118), .ZN(n660));
  XNOR2_X1  g0345(.A(n660), .B(n659), .ZN(n661));
  INV_X1    g0346(.A(81), .ZN(n662));
  MUX2_X1   g0347(.S(18), .B(349), .A(n662), .ZN(n663));
  MUX2_X1   g0348(.S(18), .B(194), .A(121), .ZN(n664));
  INV_X1    g0349(.A(n664), .ZN(n665));
  XNOR2_X1  g0350(.A(n665), .B(n663), .ZN(n666));
  INV_X1    g0351(.A(59), .ZN(n667));
  MUX2_X1   g0352(.S(18), .B(346), .A(n667), .ZN(n668));
  MUX2_X1   g0353(.S(18), .B(195), .A(94), .ZN(n669));
  XOR2_X1   g0354(.A(n669), .B(n668), .ZN(n670));
  MUX2_X1   g0355(.S(18), .B(n410), .A(78), .ZN(n671));
  MUX2_X1   g0356(.S(18), .B(196), .A(97), .ZN(n672));
  XNOR2_X1  g0357(.A(n672), .B(n671), .ZN(n673));
  OR3_X1    g0358(.A1(n673), .A2(n670), .A3(n666), .ZN(n674));
  NOR3_X1   g0359(.A1(n674), .A2(n661), .A3(n658), .ZN(n675));
  NAND2_X1  g0360(.A1(n675), .A2(n654), .ZN(n676));
  XNOR2_X1  g0361(.A(n615), .B(n614), .ZN(n677));
  OR4_X1    g0362(.A1(n613), .A2(n608), .A3(n600), .A4(n677), .ZN(n678));
  OR3_X1    g0363(.A1(n678), .A2(n594), .A3(n591), .ZN(n679));
  NOR2_X1   g0364(.A1(70), .A2(18), .ZN(n680));
  MUX2_X1   g0365(.S(18), .B(198), .A(41), .ZN(n681));
  AND2_X1   g0366(.A1(n681), .A2(n325), .ZN(n682));
  XOR2_X1   g0367(.A(n682), .B(n680), .ZN(n683));
  MUX2_X1   g0368(.S(18), .B(n458), .A(73), .ZN(n684));
  AND2_X1   g0369(.A1(204), .A2(18), .ZN(n685));
  AOI21_X1  g0370(.A(n685), .B1(103), .B2(n325), .ZN(n686));
  XOR2_X1   g0371(.A(n686), .B(n684), .ZN(n687));
  INV_X1    g0372(.A(75), .ZN(n688));
  MUX2_X1   g0373(.S(18), .B(319), .A(n688), .ZN(n689));
  MUX2_X1   g0374(.S(18), .B(205), .A(23), .ZN(n690));
  XNOR2_X1  g0375(.A(n690), .B(n689), .ZN(n691));
  INV_X1    g0376(.A(n691), .ZN(n692));
  MUX2_X1   g0377(.S(18), .B(n454), .A(76), .ZN(n693));
  MUX2_X1   g0378(.S(18), .B(206), .A(26), .ZN(n694));
  INV_X1    g0379(.A(n694), .ZN(n695));
  XNOR2_X1  g0380(.A(n695), .B(n693), .ZN(n696));
  INV_X1    g0381(.A(n696), .ZN(n697));
  MUX2_X1   g0382(.S(18), .B(n451), .A(74), .ZN(n698));
  MUX2_X1   g0383(.S(18), .B(207), .A(29), .ZN(n699));
  XNOR2_X1  g0384(.A(n699), .B(n698), .ZN(n700));
  NOR4_X1   g0385(.A1(n697), .A2(n692), .A3(n687), .A4(n700), .ZN(n701));
  INV_X1    g0386(.A(n701), .ZN(n702));
  MUX2_X1   g0387(.S(18), .B(n428), .A(56), .ZN(n703));
  MUX2_X1   g0388(.S(18), .B(200), .A(100), .ZN(n704));
  XNOR2_X1  g0389(.A(n704), .B(n703), .ZN(n705));
  MUX2_X1   g0390(.S(18), .B(n439), .A(53), .ZN(n706));
  MUX2_X1   g0391(.S(18), .B(203), .A(130), .ZN(n707));
  XNOR2_X1  g0392(.A(n707), .B(n706), .ZN(n708));
  MUX2_X1   g0393(.S(18), .B(n431), .A(55), .ZN(n709));
  MUX2_X1   g0394(.S(18), .B(201), .A(124), .ZN(n710));
  XNOR2_X1  g0395(.A(n710), .B(n709), .ZN(n711));
  MUX2_X1   g0396(.S(18), .B(n434), .A(54), .ZN(n712));
  MUX2_X1   g0397(.S(18), .B(202), .A(127), .ZN(n713));
  XNOR2_X1  g0398(.A(n713), .B(n712), .ZN(n714));
  NOR4_X1   g0399(.A1(n711), .A2(n708), .A3(n705), .A4(n714), .ZN(n715));
  NAND2_X1  g0400(.A1(n715), .A2(89), .ZN(n716));
  OR4_X1    g0401(.A1(n702), .A2(n683), .A3(n679), .A4(n716), .ZN(n717));
  NOR2_X1   g0402(.A1(n717), .A2(n676), .ZN(n718));
  AOI21_X1  g0403(.A(n331), .B1(n554), .B2(n552), .ZN(n719));
  AOI211_X1 g0404(.A(n641), .B(n719), .C1(n718), .C2(n574), .ZN(n720));
  NAND2_X1  g0405(.A1(n713), .A2(n712), .ZN(n721));
  NOR3_X1   g0406(.A1(n721), .A2(n711), .A3(n705), .ZN(n722));
  NAND2_X1  g0407(.A1(n707), .A2(n706), .ZN(n723));
  NOR4_X1   g0408(.A1(n714), .A2(n711), .A3(n705), .A4(n723), .ZN(n724));
  AND2_X1   g0409(.A1(n704), .A2(n703), .ZN(n725));
  NAND2_X1  g0410(.A1(n710), .A2(n709), .ZN(n726));
  NOR2_X1   g0411(.A1(n726), .A2(n705), .ZN(n727));
  NOR4_X1   g0412(.A1(n725), .A2(n724), .A3(n722), .A4(n727), .ZN(n728));
  NAND4_X1  g0413(.A1(n681), .A2(70), .A3(n325), .A4(n691), .ZN(n729));
  OR4_X1    g0414(.A1(n700), .A2(n697), .A3(n687), .A4(n729), .ZN(n730));
  INV_X1    g0415(.A(n687), .ZN(n731));
  NAND4_X1  g0416(.A1(n693), .A2(n691), .A3(n731), .A4(n694), .ZN(n732));
  NAND3_X1  g0417(.A1(n699), .A2(n698), .A3(n691), .ZN(n733));
  OR3_X1    g0418(.A1(n733), .A2(n697), .A3(n687), .ZN(n734));
  INV_X1    g0419(.A(n684), .ZN(n735));
  NOR2_X1   g0420(.A1(n686), .A2(n735), .ZN(n736));
  INV_X1    g0421(.A(n690), .ZN(n737));
  NOR3_X1   g0422(.A1(n737), .A2(n689), .A3(n687), .ZN(n738));
  NOR2_X1   g0423(.A1(n738), .A2(n736), .ZN(n739));
  NAND4_X1  g0424(.A1(n734), .A2(n732), .A3(n730), .A4(n739), .ZN(n740));
  NAND2_X1  g0425(.A1(n740), .A2(n715), .ZN(n741));
  AOI211_X1 g0426(.A(n679), .B(n676), .C1(n728), .C2(n741), .ZN(n742));
  NAND2_X1  g0427(.A1(n652), .A2(n651), .ZN(n743));
  NOR3_X1   g0428(.A1(n743), .A2(n650), .A3(n644), .ZN(n744));
  NAND2_X1  g0429(.A1(n646), .A2(n645), .ZN(n745));
  NOR4_X1   g0430(.A1(n653), .A2(n650), .A3(n644), .A4(n745), .ZN(n746));
  AND2_X1   g0431(.A1(n643), .A2(n642), .ZN(n747));
  NAND2_X1  g0432(.A1(n649), .A2(n648), .ZN(n748));
  NOR2_X1   g0433(.A1(n748), .A2(n644), .ZN(n749));
  NOR4_X1   g0434(.A1(n747), .A2(n746), .A3(n744), .A4(n749), .ZN(n750));
  INV_X1    g0435(.A(n666), .ZN(n751));
  NOR3_X1   g0436(.A1(n673), .A2(n670), .A3(n658), .ZN(n752));
  NAND4_X1  g0437(.A1(n751), .A2(n660), .A3(n659), .A4(n752), .ZN(n753));
  INV_X1    g0438(.A(n669), .ZN(n754));
  OR4_X1    g0439(.A1(n668), .A2(n666), .A3(n658), .A4(n754), .ZN(n755));
  INV_X1    g0440(.A(n656), .ZN(n756));
  NAND2_X1  g0441(.A1(n672), .A2(n671), .ZN(n757));
  NOR4_X1   g0442(.A1(n670), .A2(n666), .A3(n658), .A4(n757), .ZN(n758));
  NOR3_X1   g0443(.A1(n665), .A2(n663), .A3(n658), .ZN(n759));
  AOI211_X1 g0444(.A(n758), .B(n759), .C1(n657), .C2(n756), .ZN(n760));
  NAND3_X1  g0445(.A1(n760), .A2(n755), .A3(n753), .ZN(n761));
  NAND2_X1  g0446(.A1(n761), .A2(n654), .ZN(n762));
  AOI21_X1  g0447(.A(n679), .B1(n762), .B2(n750), .ZN(n763));
  OAI21_X1  g0448(.A(n574), .B1(n763), .B2(n742), .ZN(n764));
  NAND3_X1  g0449(.A1(n764), .A2(n720), .A3(n629), .ZN(10102));
  NAND2_X1  g0450(.A1(n368), .A2(n365), .ZN(n768));
  NOR4_X1   g0451(.A1(n443), .A2(n433), .A3(n430), .A4(n449), .ZN(n774));
  NAND4_X1  g0452(.A1(n504), .A2(n477), .A3(n523), .A4(n549), .ZN(10104));
  INV_X1    g0453(.A(367), .ZN(n787));
  NOR4_X1   g0454(.A1(n457), .A2(n329), .A3(n787), .A4(n463), .ZN(n788));
  OR4_X1    g0455(.A1(n463), .A2(n456), .A3(n453), .A4(n465), .ZN(n789));
  OR3_X1    g0456(.A1(n469), .A2(n463), .A3(n456), .ZN(n790));
  NAND4_X1  g0457(.A1(n789), .A2(n471), .A3(n468), .A4(n790), .ZN(n791));
  OR2_X1    g0458(.A1(n791), .A2(n788), .ZN(n792));
  XNOR2_X1  g0459(.A(n792), .B(n460), .ZN(10109));
  OR3_X1    g0460(.A1(n457), .A2(n329), .A3(n787), .ZN(n794));
  NOR3_X1   g0461(.A1(n465), .A2(n456), .A3(n453), .ZN(n795));
  NOR2_X1   g0462(.A1(n469), .A2(n456), .ZN(n796));
  AOI211_X1 g0463(.A(n795), .B(n796), .C1(n455), .C2(n454), .ZN(n797));
  NAND2_X1  g0464(.A1(n797), .A2(n794), .ZN(n798));
  XNOR2_X1  g0465(.A(n798), .B(n463), .ZN(10110));
  NOR3_X1   g0466(.A1(n453), .A2(n329), .A3(n787), .ZN(n800));
  OAI21_X1  g0467(.A(n469), .B1(n465), .B2(n453), .ZN(n801));
  OR2_X1    g0468(.A1(n801), .A2(n800), .ZN(n802));
  XNOR2_X1  g0469(.A(n802), .B(n456), .ZN(10111));
  OAI21_X1  g0470(.A(n465), .B1(n329), .B2(n787), .ZN(n804));
  XNOR2_X1  g0471(.A(n804), .B(n453), .ZN(10112));
  AND2_X1   g0472(.A1(n526), .A2(367), .ZN(n806));
  OR3_X1    g0473(.A1(n806), .A2(n474), .A3(n466), .ZN(n807));
  NOR3_X1   g0474(.A1(n443), .A2(n442), .A3(n433), .ZN(n808));
  OAI21_X1  g0475(.A(n446), .B1(n437), .B2(n433), .ZN(n809));
  OR2_X1    g0476(.A1(n809), .A2(n808), .ZN(n810));
  XNOR2_X1  g0477(.A(n810), .B(n430), .ZN(n811));
  INV_X1    g0478(.A(n430), .ZN(n812));
  NOR3_X1   g0479(.A1(n449), .A2(n443), .A3(n433), .ZN(n813));
  NOR3_X1   g0480(.A1(n809), .A2(n808), .A3(n813), .ZN(n814));
  XNOR2_X1  g0481(.A(n814), .B(n812), .ZN(n815));
  MUX2_X1   g0482(.S(n807), .B(n815), .A(n811), .ZN(10350));
  INV_X1    g0483(.A(n433), .ZN(n817));
  INV_X1    g0484(.A(n443), .ZN(n818));
  AOI21_X1  g0485(.A(n436), .B1(n818), .B2(n441), .ZN(n819));
  XNOR2_X1  g0486(.A(n819), .B(n817), .ZN(n820));
  NOR2_X1   g0487(.A1(n449), .A2(n443), .ZN(n821));
  AOI211_X1 g0488(.A(n436), .B(n821), .C1(n818), .C2(n441), .ZN(n822));
  XNOR2_X1  g0489(.A(n822), .B(n817), .ZN(n823));
  MUX2_X1   g0490(.S(n807), .B(n823), .A(n820), .ZN(10351));
  XNOR2_X1  g0491(.A(n443), .B(n441), .ZN(n825));
  NOR2_X1   g0492(.A1(n440), .A2(n439), .ZN(n826));
  XOR2_X1   g0493(.A(n826), .B(n443), .ZN(n827));
  MUX2_X1   g0494(.S(n807), .B(n827), .A(n825), .ZN(10352));
  XNOR2_X1  g0495(.A(n807), .B(n449), .ZN(10353));
  OAI21_X1  g0496(.A(n346), .B1(212), .B2(n325), .ZN(n830));
  OAI21_X1  g0497(.A(n346), .B1(211), .B2(n325), .ZN(n831));
  XNOR2_X1  g0498(.A(n831), .B(n830), .ZN(n832));
  AND3_X1   g0499(.A1(n346), .A2(n342), .A3(18), .ZN(n833));
  INV_X1    g0500(.A(n833), .ZN(n834));
  XOR2_X1   g0501(.A(n354), .B(n347), .ZN(n835));
  XNOR2_X1  g0502(.A(n351), .B(n339), .ZN(n836));
  AND3_X1   g0503(.A1(n836), .A2(n835), .A3(n834), .ZN(n837));
  NOR3_X1   g0504(.A1(n836), .A2(n835), .A3(n833), .ZN(n838));
  INV_X1    g0505(.A(n835), .ZN(n839));
  AND3_X1   g0506(.A1(n836), .A2(n839), .A3(n833), .ZN(n840));
  NOR3_X1   g0507(.A1(n836), .A2(n839), .A3(n834), .ZN(n841));
  NOR4_X1   g0508(.A1(n840), .A2(n838), .A3(n837), .A4(n841), .ZN(n842));
  XNOR2_X1  g0509(.A(n842), .B(n832), .ZN(n843));
  XNOR2_X1  g0510(.A(n404), .B(n401), .ZN(n844));
  XNOR2_X1  g0511(.A(n407), .B(n398), .ZN(n845));
  XNOR2_X1  g0512(.A(n845), .B(n844), .ZN(n846));
  MUX2_X1   g0513(.S(18), .B(227), .A(115), .ZN(n847));
  XNOR2_X1  g0514(.A(n847), .B(n414), .ZN(n848));
  XNOR2_X1  g0515(.A(n424), .B(n418), .ZN(n849));
  INV_X1    g0516(.A(n849), .ZN(n850));
  XNOR2_X1  g0517(.A(n421), .B(n411), .ZN(n851));
  INV_X1    g0518(.A(n851), .ZN(n852));
  NOR3_X1   g0519(.A1(n852), .A2(n850), .A3(n848), .ZN(n853));
  NOR3_X1   g0520(.A1(n851), .A2(n849), .A3(n848), .ZN(n854));
  INV_X1    g0521(.A(n848), .ZN(n855));
  NOR3_X1   g0522(.A1(n852), .A2(n849), .A3(n855), .ZN(n856));
  NOR3_X1   g0523(.A1(n851), .A2(n850), .A3(n855), .ZN(n857));
  NOR4_X1   g0524(.A1(n856), .A2(n854), .A3(n853), .A4(n857), .ZN(n858));
  XNOR2_X1  g0525(.A(n858), .B(n846), .ZN(n859));
  XNOR2_X1  g0526(.A(n440), .B(n435), .ZN(n860));
  XNOR2_X1  g0527(.A(n432), .B(n429), .ZN(n861));
  XNOR2_X1  g0528(.A(n861), .B(n860), .ZN(n862));
  MUX2_X1   g0529(.S(18), .B(239), .A(44), .ZN(n863));
  XNOR2_X1  g0530(.A(n863), .B(n464), .ZN(n864));
  XNOR2_X1  g0531(.A(n462), .B(n459), .ZN(n865));
  INV_X1    g0532(.A(n865), .ZN(n866));
  XNOR2_X1  g0533(.A(n455), .B(n452), .ZN(n867));
  INV_X1    g0534(.A(n867), .ZN(n868));
  NOR3_X1   g0535(.A1(n868), .A2(n866), .A3(n864), .ZN(n869));
  NOR3_X1   g0536(.A1(n867), .A2(n865), .A3(n864), .ZN(n870));
  INV_X1    g0537(.A(n864), .ZN(n871));
  NOR3_X1   g0538(.A1(n868), .A2(n865), .A3(n871), .ZN(n872));
  NOR3_X1   g0539(.A1(n867), .A2(n866), .A3(n871), .ZN(n873));
  NOR4_X1   g0540(.A1(n872), .A2(n870), .A3(n869), .A4(n873), .ZN(n874));
  XNOR2_X1  g0541(.A(n874), .B(n862), .ZN(n875));
  XNOR2_X1  g0542(.A(n367), .B(n364), .ZN(n876));
  XNOR2_X1  g0543(.A(n371), .B(n360), .ZN(n877));
  XNOR2_X1  g0544(.A(n877), .B(n876), .ZN(n878));
  XNOR2_X1  g0545(.A(n392), .B(n377), .ZN(n879));
  MUX2_X1   g0546(.S(18), .B(161), .A(141), .ZN(n880));
  XNOR2_X1  g0547(.A(n880), .B(n384), .ZN(n881));
  INV_X1    g0548(.A(n881), .ZN(n882));
  XNOR2_X1  g0549(.A(n388), .B(n381), .ZN(n883));
  AND3_X1   g0550(.A1(n883), .A2(n882), .A3(n879), .ZN(n884));
  NOR3_X1   g0551(.A1(n883), .A2(n881), .A3(n879), .ZN(n885));
  INV_X1    g0552(.A(n879), .ZN(n886));
  AND3_X1   g0553(.A1(n883), .A2(n881), .A3(n886), .ZN(n887));
  NOR3_X1   g0554(.A1(n883), .A2(n882), .A3(n886), .ZN(n888));
  NOR4_X1   g0555(.A1(n887), .A2(n885), .A3(n884), .A4(n888), .ZN(n889));
  XNOR2_X1  g0556(.A(n889), .B(n878), .ZN(n890));
  NOR4_X1   g0557(.A1(n875), .A2(n859), .A3(n843), .A4(n890), .ZN(n891));
  INV_X1    g0558(.A(n891), .ZN(10574));
  XNOR2_X1  g0559(.A(n712), .B(n706), .ZN(n893));
  XNOR2_X1  g0560(.A(n709), .B(n703), .ZN(n894));
  XNOR2_X1  g0561(.A(n894), .B(n893), .ZN(n895));
  INV_X1    g0562(.A(69), .ZN(n896));
  MUX2_X1   g0563(.S(18), .B(307), .A(n896), .ZN(n897));
  INV_X1    g0564(.A(70), .ZN(n898));
  MUX2_X1   g0565(.S(18), .B(310), .A(n898), .ZN(n899));
  XNOR2_X1  g0566(.A(n899), .B(n897), .ZN(n900));
  XOR2_X1   g0567(.A(n689), .B(n684), .ZN(n901));
  INV_X1    g0568(.A(n901), .ZN(n902));
  XNOR2_X1  g0569(.A(n698), .B(n693), .ZN(n903));
  INV_X1    g0570(.A(n903), .ZN(n904));
  NOR3_X1   g0571(.A1(n904), .A2(n902), .A3(n900), .ZN(n905));
  NOR3_X1   g0572(.A1(n903), .A2(n901), .A3(n900), .ZN(n906));
  INV_X1    g0573(.A(n900), .ZN(n907));
  NOR3_X1   g0574(.A1(n904), .A2(n901), .A3(n907), .ZN(n908));
  NOR3_X1   g0575(.A1(n903), .A2(n902), .A3(n907), .ZN(n909));
  NOR4_X1   g0576(.A1(n908), .A2(n906), .A3(n905), .A4(n909), .ZN(n910));
  XNOR2_X1  g0577(.A(n910), .B(n895), .ZN(n911));
  XNOR2_X1  g0578(.A(n587), .B(n580), .ZN(n912));
  XNOR2_X1  g0579(.A(n583), .B(n575), .ZN(n913));
  XNOR2_X1  g0580(.A(n913), .B(n912), .ZN(n914));
  INV_X1    g0581(.A(82), .ZN(n915));
  MUX2_X1   g0582(.S(18), .B(274), .A(n915), .ZN(n916));
  XOR2_X1   g0583(.A(n916), .B(n614), .ZN(n917));
  XNOR2_X1  g0584(.A(n595), .B(n592), .ZN(n918));
  INV_X1    g0585(.A(n918), .ZN(n919));
  XNOR2_X1  g0586(.A(n610), .B(n602), .ZN(n920));
  INV_X1    g0587(.A(n920), .ZN(n921));
  NOR3_X1   g0588(.A1(n921), .A2(n919), .A3(n917), .ZN(n922));
  NOR3_X1   g0589(.A1(n920), .A2(n918), .A3(n917), .ZN(n923));
  INV_X1    g0590(.A(n917), .ZN(n924));
  NOR3_X1   g0591(.A1(n921), .A2(n918), .A3(n924), .ZN(n925));
  NOR3_X1   g0592(.A1(n920), .A2(n919), .A3(n924), .ZN(n926));
  NOR4_X1   g0593(.A1(n925), .A2(n923), .A3(n922), .A4(n926), .ZN(n927));
  XNOR2_X1  g0594(.A(n927), .B(n914), .ZN(n928));
  XNOR2_X1  g0595(.A(n651), .B(n645), .ZN(n929));
  XNOR2_X1  g0596(.A(n648), .B(n642), .ZN(n930));
  XNOR2_X1  g0597(.A(n930), .B(n929), .ZN(n931));
  INV_X1    g0598(.A(58), .ZN(n932));
  MUX2_X1   g0599(.S(18), .B(337), .A(n932), .ZN(n933));
  XOR2_X1   g0600(.A(n933), .B(n659), .ZN(n934));
  XNOR2_X1  g0601(.A(n663), .B(n656), .ZN(n935));
  INV_X1    g0602(.A(n935), .ZN(n936));
  XOR2_X1   g0603(.A(n671), .B(n668), .ZN(n937));
  INV_X1    g0604(.A(n937), .ZN(n938));
  NOR3_X1   g0605(.A1(n938), .A2(n936), .A3(n934), .ZN(n939));
  NOR3_X1   g0606(.A1(n937), .A2(n935), .A3(n934), .ZN(n940));
  INV_X1    g0607(.A(n934), .ZN(n941));
  NOR3_X1   g0608(.A1(n938), .A2(n935), .A3(n941), .ZN(n942));
  NOR3_X1   g0609(.A1(n937), .A2(n936), .A3(n941), .ZN(n943));
  NOR4_X1   g0610(.A1(n942), .A2(n940), .A3(n939), .A4(n943), .ZN(n944));
  XNOR2_X1  g0611(.A(n944), .B(n931), .ZN(n945));
  INV_X1    g0612(.A(245), .ZN(n946));
  MUX2_X1   g0613(.S(18), .B(263), .A(n946), .ZN(n947));
  INV_X1    g0614(.A(271), .ZN(n948));
  MUX2_X1   g0615(.S(n325), .B(n948), .A(267), .ZN(n949));
  XNOR2_X1  g0616(.A(n949), .B(n947), .ZN(n950));
  INV_X1    g0617(.A(114), .ZN(n951));
  MUX2_X1   g0618(.S(18), .B(248), .A(n951), .ZN(n952));
  XOR2_X1   g0619(.A(n952), .B(n561), .ZN(n953));
  XOR2_X1   g0620(.A(n563), .B(n557), .ZN(n954));
  INV_X1    g0621(.A(n954), .ZN(n955));
  XNOR2_X1  g0622(.A(n569), .B(n566), .ZN(n956));
  INV_X1    g0623(.A(n956), .ZN(n957));
  NOR3_X1   g0624(.A1(n957), .A2(n955), .A3(n953), .ZN(n958));
  NOR3_X1   g0625(.A1(n956), .A2(n954), .A3(n953), .ZN(n959));
  INV_X1    g0626(.A(n953), .ZN(n960));
  NOR3_X1   g0627(.A1(n957), .A2(n954), .A3(n960), .ZN(n961));
  NOR3_X1   g0628(.A1(n956), .A2(n955), .A3(n960), .ZN(n962));
  NOR4_X1   g0629(.A1(n961), .A2(n959), .A3(n958), .A4(n962), .ZN(n963));
  XNOR2_X1  g0630(.A(n963), .B(n950), .ZN(n964));
  NOR4_X1   g0631(.A1(n945), .A2(n928), .A3(n911), .A4(n964), .ZN(n965));
  INV_X1    g0632(.A(n965), .ZN(10575));
  OAI21_X1  g0633(.A(n346), .B1(165), .B2(n325), .ZN(n967));
  OAI21_X1  g0634(.A(n346), .B1(164), .B2(n325), .ZN(n968));
  XNOR2_X1  g0635(.A(n968), .B(n967), .ZN(n969));
  NAND2_X1  g0636(.A1(170), .A2(18), .ZN(n970));
  AND3_X1   g0637(.A1(n970), .A2(n346), .A3(18), .ZN(n971));
  INV_X1    g0638(.A(n971), .ZN(n972));
  XNOR2_X1  g0639(.A(n564), .B(n558), .ZN(n973));
  XNOR2_X1  g0640(.A(n570), .B(n567), .ZN(n974));
  AND3_X1   g0641(.A1(n974), .A2(n973), .A3(n972), .ZN(n975));
  NOR3_X1   g0642(.A1(n974), .A2(n973), .A3(n971), .ZN(n976));
  INV_X1    g0643(.A(n973), .ZN(n977));
  AND3_X1   g0644(.A1(n974), .A2(n977), .A3(n971), .ZN(n978));
  NOR3_X1   g0645(.A1(n974), .A2(n977), .A3(n972), .ZN(n979));
  NOR4_X1   g0646(.A1(n978), .A2(n976), .A3(n975), .A4(n979), .ZN(n980));
  XNOR2_X1  g0647(.A(n980), .B(n969), .ZN(n981));
  XNOR2_X1  g0648(.A(n652), .B(n646), .ZN(n982));
  XNOR2_X1  g0649(.A(n649), .B(n643), .ZN(n983));
  XNOR2_X1  g0650(.A(n983), .B(n982), .ZN(n984));
  MUX2_X1   g0651(.S(18), .B(197), .A(115), .ZN(n985));
  XNOR2_X1  g0652(.A(n985), .B(n660), .ZN(n986));
  XNOR2_X1  g0653(.A(n664), .B(n657), .ZN(n987));
  INV_X1    g0654(.A(n987), .ZN(n988));
  XNOR2_X1  g0655(.A(n672), .B(n669), .ZN(n989));
  INV_X1    g0656(.A(n989), .ZN(n990));
  NOR3_X1   g0657(.A1(n990), .A2(n988), .A3(n986), .ZN(n991));
  NOR3_X1   g0658(.A1(n989), .A2(n987), .A3(n986), .ZN(n992));
  INV_X1    g0659(.A(n986), .ZN(n993));
  NOR3_X1   g0660(.A1(n990), .A2(n987), .A3(n993), .ZN(n994));
  NOR3_X1   g0661(.A1(n989), .A2(n988), .A3(n993), .ZN(n995));
  NOR4_X1   g0662(.A1(n994), .A2(n992), .A3(n991), .A4(n995), .ZN(n996));
  XNOR2_X1  g0663(.A(n996), .B(n984), .ZN(n997));
  XNOR2_X1  g0664(.A(n713), .B(n707), .ZN(n998));
  XNOR2_X1  g0665(.A(n710), .B(n704), .ZN(n999));
  XNOR2_X1  g0666(.A(n999), .B(n998), .ZN(n1000));
  MUX2_X1   g0667(.S(18), .B(208), .A(44), .ZN(n1001));
  XNOR2_X1  g0668(.A(n1001), .B(n681), .ZN(n1002));
  INV_X1    g0669(.A(n1002), .ZN(n1003));
  XNOR2_X1  g0670(.A(n737), .B(n686), .ZN(n1004));
  XNOR2_X1  g0671(.A(n699), .B(n694), .ZN(n1005));
  AND3_X1   g0672(.A1(n1005), .A2(n1004), .A3(n1003), .ZN(n1006));
  NOR3_X1   g0673(.A1(n1005), .A2(n1004), .A3(n1002), .ZN(n1007));
  INV_X1    g0674(.A(n1004), .ZN(n1008));
  AND3_X1   g0675(.A1(n1005), .A2(n1008), .A3(n1002), .ZN(n1009));
  NOR3_X1   g0676(.A1(n1005), .A2(n1008), .A3(n1003), .ZN(n1010));
  NOR4_X1   g0677(.A1(n1009), .A2(n1007), .A3(n1006), .A4(n1010), .ZN(n1011));
  XNOR2_X1  g0678(.A(n1011), .B(n1000), .ZN(n1012));
  XOR2_X1   g0679(.A(n589), .B(n581), .ZN(n1013));
  XOR2_X1   g0680(.A(n584), .B(n577), .ZN(n1014));
  XNOR2_X1  g0681(.A(n1014), .B(n1013), .ZN(n1015));
  XNOR2_X1  g0682(.A(n598), .B(n593), .ZN(n1016));
  MUX2_X1   g0683(.S(18), .B(181), .A(141), .ZN(n1017));
  XNOR2_X1  g0684(.A(n1017), .B(n615), .ZN(n1018));
  INV_X1    g0685(.A(n1018), .ZN(n1019));
  XNOR2_X1  g0686(.A(n611), .B(n603), .ZN(n1020));
  AND3_X1   g0687(.A1(n1020), .A2(n1019), .A3(n1016), .ZN(n1021));
  NOR3_X1   g0688(.A1(n1020), .A2(n1018), .A3(n1016), .ZN(n1022));
  INV_X1    g0689(.A(n1016), .ZN(n1023));
  AND3_X1   g0690(.A1(n1020), .A2(n1018), .A3(n1023), .ZN(n1024));
  NOR3_X1   g0691(.A1(n1020), .A2(n1019), .A3(n1023), .ZN(n1025));
  NOR4_X1   g0692(.A1(n1024), .A2(n1022), .A3(n1021), .A4(n1025), .ZN(n1026));
  XNOR2_X1  g0693(.A(n1026), .B(n1015), .ZN(n1027));
  NOR4_X1   g0694(.A1(n1012), .A2(n997), .A3(n981), .A4(n1027), .ZN(n1028));
  INV_X1    g0695(.A(n1028), .ZN(10576));
  OAI211_X1 g0696(.A(n331), .B(382), .C1(n948), .C2(n946), .ZN(n1030));
  NOR4_X1   g0697(.A1(n742), .A2(n718), .A3(n628), .A4(n763), .ZN(n1031));
  OAI21_X1  g0698(.A(n640), .B1(n1031), .B2(n573), .ZN(n1032));
  MUX2_X1   g0699(.S(n1032), .B(n1030), .A(n719), .ZN(10628));
  NAND2_X1  g0700(.A1(n476), .A2(n427), .ZN(n1034));
  AND2_X1   g0701(.A1(n527), .A2(n502), .ZN(n1035));
  NAND2_X1  g0702(.A1(n1035), .A2(n1034), .ZN(n1036));
  XNOR2_X1  g0703(.A(n1036), .B(n385), .ZN(10632));
  AND3_X1   g0704(.A1(n476), .A2(n427), .A3(n396), .ZN(n1038));
  NOR4_X1   g0705(.A1(n528), .A2(n503), .A3(n1038), .A4(n548), .ZN(n1039));
  XOR2_X1   g0706(.A(n1039), .B(n344), .ZN(10641));
  INV_X1    g0707(.A(n654), .ZN(n1041));
  INV_X1    g0708(.A(n715), .ZN(n1042));
  NOR2_X1   g0709(.A1(n702), .A2(n683), .ZN(n1043));
  AOI21_X1  g0710(.A(n740), .B1(n1043), .B2(89), .ZN(n1044));
  OAI21_X1  g0711(.A(n728), .B1(n1044), .B2(n1042), .ZN(n1045));
  AOI21_X1  g0712(.A(n761), .B1(n1045), .B2(n675), .ZN(n1046));
  OAI21_X1  g0713(.A(n750), .B1(n1046), .B2(n1041), .ZN(10704));
  NOR2_X1   g0714(.A1(n505), .A2(n336), .ZN(n1048));
  INV_X1    g0715(.A(n1048), .ZN(n1049));
  INV_X1    g0716(.A(n356), .ZN(n1050));
  OAI21_X1  g0717(.A(n521), .B1(n1039), .B2(n1050), .ZN(n1053));
  MUX2_X1   g0718(.S(n1053), .B(n1049), .A(n505), .ZN(10706));
  AOI21_X1  g0719(.A(n385), .B1(n1035), .B2(n1034), .ZN(n1055));
  AND2_X1   g0720(.A1(n1055), .A2(n542), .ZN(n1056));
  AND3_X1   g0721(.A1(n394), .A2(n388), .A3(n387), .ZN(n1057));
  AND3_X1   g0722(.A1(n543), .A2(n542), .A3(n394), .ZN(n1058));
  NOR3_X1   g0723(.A1(n545), .A2(n393), .A3(n389), .ZN(n1059));
  OR4_X1    g0724(.A1(n1058), .A2(n1057), .A3(n537), .A4(n1059), .ZN(n1060));
  AOI21_X1  g0725(.A(n1060), .B1(n1056), .B2(n394), .ZN(n1061));
  XOR2_X1   g0726(.A(n1061), .B(n378), .ZN(10711));
  NOR2_X1   g0727(.A1(n545), .A2(n389), .ZN(n1063));
  AOI221_X1 g0728(.A(n1063), .B1(n542), .B2(n543), .C1(n388), .C2(n387), .ZN(n1064));
  INV_X1    g0729(.A(n1064), .ZN(n1065));
  AOI21_X1  g0730(.A(n1065), .B1(n1055), .B2(n542), .ZN(n1066));
  XNOR2_X1  g0731(.A(n1066), .B(n394), .ZN(10712));
  INV_X1    g0732(.A(n382), .ZN(n1068));
  INV_X1    g0733(.A(n543), .ZN(n1069));
  OAI21_X1  g0734(.A(n545), .B1(n1069), .B2(n382), .ZN(n1070));
  AOI21_X1  g0735(.A(n1070), .B1(n1055), .B2(n1068), .ZN(n1071));
  XOR2_X1   g0736(.A(n1071), .B(n389), .ZN(10713));
  NOR2_X1   g0737(.A1(n1055), .A2(n543), .ZN(n1073));
  XNOR2_X1  g0738(.A(n1073), .B(n1068), .ZN(10714));
  NOR4_X1   g0739(.A1(n507), .A2(n344), .A3(n340), .A4(n1039), .ZN(n1075));
  NOR2_X1   g0740(.A1(n513), .A2(n512), .ZN(n1076));
  XNOR2_X1  g0741(.A(n339), .B(254), .ZN(n1077));
  AND4_X1   g0742(.A1(n355), .A2(n352), .A3(n1077), .A4(n509), .ZN(n1078));
  NOR3_X1   g0743(.A1(n515), .A2(n512), .A3(n507), .ZN(n1079));
  OR4_X1    g0744(.A1(n1078), .A2(n518), .A3(n1076), .A4(n1079), .ZN(n1080));
  AOI21_X1  g0745(.A(n1080), .B1(n1075), .B2(n355), .ZN(n1081));
  XOR2_X1   g0746(.A(n1081), .B(n348), .ZN(10715));
  NAND3_X1  g0747(.A1(n509), .A2(n352), .A3(n1077), .ZN(n1083));
  OR2_X1    g0748(.A1(n515), .A2(n507), .ZN(n1084));
  AND3_X1   g0749(.A1(n1084), .A2(n1083), .A3(n513), .ZN(n1085));
  INV_X1    g0750(.A(n1085), .ZN(n1086));
  NOR2_X1   g0751(.A1(n1086), .A2(n1075), .ZN(n1087));
  XNOR2_X1  g0752(.A(n1087), .B(n355), .ZN(10716));
  NOR3_X1   g0753(.A1(n1039), .A2(n344), .A3(n340), .ZN(n1089));
  INV_X1    g0754(.A(n509), .ZN(n1090));
  OAI21_X1  g0755(.A(n515), .B1(n1090), .B2(n340), .ZN(n1091));
  NOR2_X1   g0756(.A1(n1091), .A2(n1089), .ZN(n1092));
  XOR2_X1   g0757(.A(n1092), .B(n507), .ZN(10717));
  OAI21_X1  g0758(.A(n1090), .B1(n1039), .B2(n344), .ZN(n1094));
  XNOR2_X1  g0759(.A(n1094), .B(n340), .ZN(10718));
  NOR4_X1   g0760(.A1(884), .A2(883), .A3(882), .A4(885), .ZN(n1096));
  NAND4_X1  g0761(.A1(n1028), .A2(n965), .A3(n891), .A4(n1096), .ZN(10729));
  MUX2_X1   g0762(.S(n1053), .B(n1049), .A(n505), .ZN(10759));
  INV_X1    g0763(.A(n547), .ZN(n1101));
  AOI21_X1  g0764(.A(n395), .B1(n1035), .B2(n1034), .ZN(n1102));
  OR2_X1    g0765(.A1(n1102), .A2(n1101), .ZN(n1103));
  AND2_X1   g0766(.A1(n529), .A2(n373), .ZN(n1104));
  INV_X1    g0767(.A(n368), .ZN(n1105));
  INV_X1    g0768(.A(n531), .ZN(n1106));
  NOR3_X1   g0769(.A1(n1106), .A2(n372), .A3(n1105), .ZN(n1107));
  NOR3_X1   g0770(.A1(n1107), .A2(n534), .A3(n1104), .ZN(n1108));
  XNOR2_X1  g0771(.A(n1108), .B(n362), .ZN(n1109));
  NOR2_X1   g0772(.A1(n768), .A2(n372), .ZN(n1110));
  NOR4_X1   g0773(.A1(n1110), .A2(n534), .A3(n1104), .A4(n1107), .ZN(n1111));
  XNOR2_X1  g0774(.A(n1111), .B(n362), .ZN(n1112));
  MUX2_X1   g0775(.S(n1103), .B(n1112), .A(n1109), .ZN(10760));
  AOI21_X1  g0776(.A(n529), .B1(n531), .B2(n368), .ZN(n1114));
  XNOR2_X1  g0777(.A(n1114), .B(n373), .ZN(n1115));
  AND2_X1   g0778(.A1(n1114), .A2(n768), .ZN(n1116));
  XNOR2_X1  g0779(.A(n1116), .B(n373), .ZN(n1117));
  MUX2_X1   g0780(.S(n1103), .B(n1117), .A(n1115), .ZN(10761));
  XNOR2_X1  g0781(.A(n1106), .B(n368), .ZN(n1119));
  NOR2_X1   g0782(.A1(n364), .A2(n579), .ZN(n1120));
  XNOR2_X1  g0783(.A(n1120), .B(n368), .ZN(n1121));
  MUX2_X1   g0784(.S(n1103), .B(n1121), .A(n1119), .ZN(10762));
  INV_X1    g0785(.A(n365), .ZN(n1123));
  XNOR2_X1  g0786(.A(n1103), .B(n1123), .ZN(10763));
  INV_X1    g0787(.A(n448), .ZN(n1125));
  AOI21_X1  g0788(.A(n1125), .B1(n807), .B2(n774), .ZN(n1126));
  XOR2_X1   g0789(.A(n1126), .B(n415), .ZN(10827));
  NOR2_X1   g0790(.A1(n334), .A2(n331), .ZN(n1128));
  XNOR2_X1  g0791(.A(n1128), .B(n333), .ZN(n1129));
  NAND2_X1  g0792(.A1(n334), .A2(n331), .ZN(n1130));
  XNOR2_X1  g0793(.A(n1130), .B(n333), .ZN(n1131));
  MUX2_X1   g0794(.S(n1053), .B(n1131), .A(n1129), .ZN(10837));
  XNOR2_X1  g0795(.A(n1053), .B(n335), .ZN(10839));
  INV_X1    g0796(.A(n492), .ZN(n1134));
  NOR4_X1   g0797(.A1(n1134), .A2(n425), .A3(n415), .A4(n1126), .ZN(n1135));
  AND3_X1   g0798(.A1(n491), .A2(n421), .A3(n420), .ZN(n1136));
  AND3_X1   g0799(.A1(n493), .A2(n492), .A3(n491), .ZN(n1137));
  NOR3_X1   g0800(.A1(n496), .A2(n425), .A3(n422), .ZN(n1138));
  OR4_X1    g0801(.A1(n1137), .A2(n499), .A3(n1136), .A4(n1138), .ZN(n1139));
  NOR2_X1   g0802(.A1(n1139), .A2(n1135), .ZN(n1140));
  XNOR2_X1  g0803(.A(n1140), .B(n490), .ZN(10868));
  OR3_X1    g0804(.A1(n1126), .A2(n1134), .A3(n415), .ZN(n1142));
  NOR2_X1   g0805(.A1(n496), .A2(n422), .ZN(n1143));
  AOI221_X1 g0806(.A(n1143), .B1(n492), .B2(n493), .C1(n421), .C2(n420), .ZN(n1144));
  AND2_X1   g0807(.A1(n1144), .A2(n1142), .ZN(n1145));
  XNOR2_X1  g0808(.A(n1145), .B(n491), .ZN(10869));
  NOR3_X1   g0809(.A1(n1126), .A2(n415), .A3(n412), .ZN(n1147));
  INV_X1    g0810(.A(n493), .ZN(n1148));
  OAI21_X1  g0811(.A(n496), .B1(n1148), .B2(n412), .ZN(n1149));
  OR2_X1    g0812(.A1(n1149), .A2(n1147), .ZN(n1150));
  XNOR2_X1  g0813(.A(n1150), .B(n422), .ZN(10870));
  OAI21_X1  g0814(.A(n1148), .B1(n1126), .B2(n415), .ZN(n1152));
  XNOR2_X1  g0815(.A(n1152), .B(n412), .ZN(10871));
  AOI21_X1  g0816(.A(n501), .B1(n1264), .B2(n426), .ZN(n1155));
  NOR2_X1   g0817(.A1(n479), .A2(n408), .ZN(n1156));
  AND3_X1   g0818(.A1(n484), .A2(n483), .A3(n482), .ZN(n1157));
  OR3_X1    g0819(.A1(n1157), .A2(n487), .A3(n1156), .ZN(n1158));
  XNOR2_X1  g0820(.A(n1158), .B(n399), .ZN(n1159));
  NOR3_X1   g0821(.A1(n408), .A2(n405), .A3(n402), .ZN(n1160));
  NOR4_X1   g0822(.A1(n1160), .A2(n487), .A3(n1156), .A4(n1157), .ZN(n1161));
  XNOR2_X1  g0823(.A(n1161), .B(n481), .ZN(n1162));
  MUX2_X1   g0824(.S(n1155), .B(n1159), .A(n1162), .ZN(10905));
  AOI21_X1  g0825(.A(n478), .B1(n484), .B2(n482), .ZN(n1164));
  XNOR2_X1  g0826(.A(n1164), .B(n483), .ZN(n1165));
  NOR2_X1   g0827(.A1(n405), .A2(n402), .ZN(n1166));
  AOI211_X1 g0828(.A(n478), .B(n1166), .C1(n484), .C2(n482), .ZN(n1167));
  XNOR2_X1  g0829(.A(n1167), .B(n483), .ZN(n1168));
  MUX2_X1   g0830(.S(n1155), .B(n1165), .A(n1168), .ZN(10906));
  XNOR2_X1  g0831(.A(n484), .B(n405), .ZN(n1170));
  NOR2_X1   g0832(.A1(n401), .A2(n400), .ZN(n1171));
  XOR2_X1   g0833(.A(n1171), .B(n405), .ZN(n1172));
  MUX2_X1   g0834(.S(n1155), .B(n1170), .A(n1172), .ZN(10907));
  XOR2_X1   g0835(.A(n1155), .B(n402), .ZN(10908));
  XNOR2_X1  g0836(.A(n1064), .B(n543), .ZN(n1175));
  XNOR2_X1  g0837(.A(n1175), .B(n1070), .ZN(n1176));
  XNOR2_X1  g0838(.A(n1176), .B(n1060), .ZN(n1177));
  XNOR2_X1  g0839(.A(n1177), .B(n385), .ZN(n1178));
  XNOR2_X1  g0840(.A(n1178), .B(n382), .ZN(n1179));
  XNOR2_X1  g0841(.A(n1179), .B(n378), .ZN(n1180));
  XNOR2_X1  g0842(.A(n1180), .B(n389), .ZN(n1181));
  OR2_X1    g0843(.A1(n1181), .A2(n394), .ZN(n1182));
  AND3_X1   g0844(.A1(n527), .A2(n502), .A3(n1034), .ZN(n1185));
  AOI21_X1  g0845(.A(n1036), .B1(n1181), .B2(n394), .ZN(n1187));
  NOR4_X1   g0846(.A1(n389), .A2(n385), .A3(n382), .A4(n393), .ZN(n1188));
  NOR2_X1   g0847(.A1(n1188), .A2(n1060), .ZN(n1189));
  NOR2_X1   g0848(.A1(n1070), .A2(n386), .ZN(n1190));
  OR3_X1    g0849(.A1(n389), .A2(n385), .A3(n382), .ZN(n1191));
  NAND2_X1  g0850(.A1(n1191), .A2(n1064), .ZN(n1192));
  NOR2_X1   g0851(.A1(n384), .A2(n383), .ZN(n1193));
  XNOR2_X1  g0852(.A(n1193), .B(n1192), .ZN(n1194));
  XNOR2_X1  g0853(.A(n1194), .B(n1190), .ZN(n1195));
  XNOR2_X1  g0854(.A(n1195), .B(n1189), .ZN(n1196));
  XNOR2_X1  g0855(.A(n1196), .B(n385), .ZN(n1197));
  XNOR2_X1  g0856(.A(n1197), .B(n382), .ZN(n1198));
  XNOR2_X1  g0857(.A(n1198), .B(n378), .ZN(n1199));
  XNOR2_X1  g0858(.A(n1199), .B(n389), .ZN(n1200));
  XNOR2_X1  g0859(.A(n1200), .B(n394), .ZN(n1201));
  AOI22_X1  g0860(.A1(n1187), .A2(n1182), .B1(n1036), .B2(n1201), .ZN(n1202));
  XOR2_X1   g0861(.A(n1120), .B(n1116), .ZN(n1203));
  XNOR2_X1  g0862(.A(n1203), .B(n1111), .ZN(n1204));
  XNOR2_X1  g0863(.A(n1204), .B(n1123), .ZN(n1205));
  XNOR2_X1  g0864(.A(n1205), .B(n1105), .ZN(n1206));
  XNOR2_X1  g0865(.A(n1206), .B(n361), .ZN(n1207));
  XNOR2_X1  g0866(.A(n1207), .B(n372), .ZN(n1208));
  NOR3_X1   g0867(.A1(n1208), .A2(n1036), .A3(n547), .ZN(n1209));
  AOI211_X1 g0868(.A(n1185), .B(n1208), .C1(n547), .C2(n395), .ZN(n1210));
  INV_X1    g0869(.A(n395), .ZN(n1211));
  XNOR2_X1  g0870(.A(n1114), .B(n1106), .ZN(n1212));
  XNOR2_X1  g0871(.A(n1212), .B(n1108), .ZN(n1213));
  XNOR2_X1  g0872(.A(n1213), .B(n1123), .ZN(n1214));
  XNOR2_X1  g0873(.A(n1214), .B(n1105), .ZN(n1215));
  XNOR2_X1  g0874(.A(n1215), .B(n361), .ZN(n1216));
  XNOR2_X1  g0875(.A(n1216), .B(n372), .ZN(n1217));
  AOI211_X1 g0876(.A(n1101), .B(n1217), .C1(n1036), .C2(n1211), .ZN(n1218));
  NOR3_X1   g0877(.A1(n1218), .A2(n1210), .A3(n1209), .ZN(n1219));
  XNOR2_X1  g0878(.A(n1219), .B(n1202), .ZN(11333));
  INV_X1    g0879(.A(n1039), .ZN(n1221));
  XNOR2_X1  g0880(.A(n1085), .B(n509), .ZN(n1222));
  XNOR2_X1  g0881(.A(n1222), .B(n1091), .ZN(n1223));
  XNOR2_X1  g0882(.A(n1223), .B(n1080), .ZN(n1224));
  XNOR2_X1  g0883(.A(n1224), .B(n344), .ZN(n1225));
  XNOR2_X1  g0884(.A(n1225), .B(n340), .ZN(n1226));
  XNOR2_X1  g0885(.A(n1226), .B(n348), .ZN(n1227));
  XNOR2_X1  g0886(.A(n1227), .B(n352), .ZN(n1228));
  OR2_X1    g0887(.A1(n1228), .A2(n512), .ZN(n1229));
  AOI21_X1  g0888(.A(n1221), .B1(n1228), .B2(n512), .ZN(n1230));
  NOR4_X1   g0889(.A1(n507), .A2(n344), .A3(n340), .A4(n512), .ZN(n1231));
  NOR2_X1   g0890(.A1(n1231), .A2(n1080), .ZN(n1232));
  NOR2_X1   g0891(.A1(n1091), .A2(n345), .ZN(n1233));
  OR3_X1    g0892(.A1(n507), .A2(n344), .A3(n340), .ZN(n1234));
  NAND4_X1  g0893(.A1(n1084), .A2(n1083), .A3(n513), .A4(n1234), .ZN(n1235));
  NOR2_X1   g0894(.A1(n343), .A2(n341), .ZN(n1236));
  XNOR2_X1  g0895(.A(n1236), .B(n1235), .ZN(n1237));
  XNOR2_X1  g0896(.A(n1237), .B(n1233), .ZN(n1238));
  XNOR2_X1  g0897(.A(n1238), .B(n1232), .ZN(n1239));
  XNOR2_X1  g0898(.A(n1239), .B(n344), .ZN(n1240));
  XNOR2_X1  g0899(.A(n1240), .B(n340), .ZN(n1241));
  XNOR2_X1  g0900(.A(n1241), .B(n348), .ZN(n1242));
  XNOR2_X1  g0901(.A(n1242), .B(n507), .ZN(n1243));
  XNOR2_X1  g0902(.A(n1243), .B(n355), .ZN(n1244));
  AOI22_X1  g0903(.A1(n1230), .A2(n1229), .B1(n1221), .B2(n1244), .ZN(n1245));
  NOR3_X1   g0904(.A1(n1129), .A2(n1221), .A3(n521), .ZN(n1248));
  AOI211_X1 g0905(.A(n1039), .B(n1129), .C1(n1050), .C2(n521), .ZN(n1249));
  AND3_X1   g0906(.A1(382), .A2(263), .A3(n331), .ZN(n1250));
  XNOR2_X1  g0907(.A(n1250), .B(n333), .ZN(n1251));
  AOI211_X1 g0908(.A(n522), .B(n1251), .C1(n1221), .C2(n356), .ZN(n1252));
  NOR3_X1   g0909(.A1(n1252), .A2(n1249), .A3(n1248), .ZN(n1253));
  XNOR2_X1  g0910(.A(n1253), .B(n1245), .ZN(11334));
  XNOR2_X1  g0911(.A(n1144), .B(n493), .ZN(n1255));
  XNOR2_X1  g0912(.A(n1255), .B(n1149), .ZN(n1256));
  XNOR2_X1  g0913(.A(n1256), .B(n1139), .ZN(n1257));
  XNOR2_X1  g0914(.A(n1257), .B(n415), .ZN(n1258));
  XNOR2_X1  g0915(.A(n1258), .B(n412), .ZN(n1259));
  XNOR2_X1  g0916(.A(n1259), .B(n419), .ZN(n1260));
  XNOR2_X1  g0917(.A(n1260), .B(n422), .ZN(n1261));
  OR2_X1    g0918(.A1(n1261), .A2(n491), .ZN(n1262));
  AOI211_X1 g0919(.A(n474), .B(n466), .C1(367), .C2(n526), .ZN(n1263));
  OAI21_X1  g0920(.A(n448), .B1(n1263), .B2(n450), .ZN(n1264));
  AOI21_X1  g0921(.A(n1264), .B1(n1261), .B2(n491), .ZN(n1265));
  NOR4_X1   g0922(.A1(n422), .A2(n415), .A3(n412), .A4(n425), .ZN(n1266));
  NOR2_X1   g0923(.A1(n1266), .A2(n1139), .ZN(n1267));
  OAI211_X1 g0924(.A(n416), .B(n496), .C1(n1148), .C2(n412), .ZN(n1268));
  OR3_X1    g0925(.A1(n422), .A2(n415), .A3(n412), .ZN(n1269));
  NAND2_X1  g0926(.A1(n1269), .A2(n1144), .ZN(n1270));
  NOR2_X1   g0927(.A1(n414), .A2(n413), .ZN(n1271));
  XOR2_X1   g0928(.A(n1271), .B(n1270), .ZN(n1272));
  XNOR2_X1  g0929(.A(n1272), .B(n1268), .ZN(n1273));
  XNOR2_X1  g0930(.A(n1273), .B(n1267), .ZN(n1274));
  XNOR2_X1  g0931(.A(n1274), .B(n415), .ZN(n1275));
  XNOR2_X1  g0932(.A(n1275), .B(n412), .ZN(n1276));
  XNOR2_X1  g0933(.A(n1276), .B(n419), .ZN(n1277));
  XNOR2_X1  g0934(.A(n1277), .B(n422), .ZN(n1278));
  XNOR2_X1  g0935(.A(n1278), .B(n491), .ZN(n1279));
  AOI22_X1  g0936(.A1(n1265), .A2(n1262), .B1(n1264), .B2(n1279), .ZN(n1280));
  XOR2_X1   g0937(.A(n1171), .B(n1167), .ZN(n1281));
  XNOR2_X1  g0938(.A(n1281), .B(n1161), .ZN(n1282));
  XNOR2_X1  g0939(.A(n1282), .B(n402), .ZN(n1283));
  XNOR2_X1  g0940(.A(n1283), .B(n405), .ZN(n1284));
  XNOR2_X1  g0941(.A(n1284), .B(n399), .ZN(n1285));
  XNOR2_X1  g0942(.A(n1285), .B(n408), .ZN(n1286));
  OAI211_X1 g0943(.A(n501), .B(n448), .C1(n450), .C2(n1263), .ZN(n1287));
  NOR2_X1   g0944(.A1(n1287), .A2(n1286), .ZN(n1288));
  OAI21_X1  g0945(.A(n1264), .B1(n426), .B2(n501), .ZN(n1289));
  NOR2_X1   g0946(.A1(n1289), .A2(n1286), .ZN(n1290));
  XNOR2_X1  g0947(.A(n1164), .B(n484), .ZN(n1291));
  XNOR2_X1  g0948(.A(n1291), .B(n1158), .ZN(n1292));
  XNOR2_X1  g0949(.A(n1292), .B(n402), .ZN(n1293));
  XNOR2_X1  g0950(.A(n1293), .B(n405), .ZN(n1294));
  XNOR2_X1  g0951(.A(n1294), .B(n399), .ZN(n1295));
  XNOR2_X1  g0952(.A(n1295), .B(n408), .ZN(n1296));
  AOI211_X1 g0953(.A(n501), .B(n1296), .C1(n1264), .C2(n426), .ZN(n1297));
  NOR3_X1   g0954(.A1(n1297), .A2(n1290), .A3(n1288), .ZN(n1298));
  XNOR2_X1  g0955(.A(n1298), .B(n1280), .ZN(11340));
  XOR2_X1   g0956(.A(n797), .B(n465), .ZN(n1300));
  XNOR2_X1  g0957(.A(n1300), .B(n801), .ZN(n1301));
  XNOR2_X1  g0958(.A(n1301), .B(n791), .ZN(n1302));
  XNOR2_X1  g0959(.A(n1302), .B(n329), .ZN(n1303));
  XNOR2_X1  g0960(.A(n1303), .B(n453), .ZN(n1304));
  XNOR2_X1  g0961(.A(n1304), .B(n460), .ZN(n1305));
  XOR2_X1   g0962(.A(n1305), .B(n456), .ZN(n1306));
  OR2_X1    g0963(.A1(n1306), .A2(n463), .ZN(n1307));
  AOI21_X1  g0964(.A(367), .B1(n1306), .B2(n463), .ZN(n1308));
  NOR4_X1   g0965(.A1(n456), .A2(n453), .A3(n329), .A4(n463), .ZN(n1309));
  NOR2_X1   g0966(.A1(n1309), .A2(n791), .ZN(n1310));
  NOR2_X1   g0967(.A1(n453), .A2(n329), .ZN(n1311));
  NOR2_X1   g0968(.A1(n801), .A2(n1311), .ZN(n1312));
  OR3_X1    g0969(.A1(n456), .A2(n453), .A3(n329), .ZN(n1313));
  NAND2_X1  g0970(.A1(n1313), .A2(n797), .ZN(n1314));
  NOR3_X1   g0971(.A1(n464), .A2(n327), .A3(18), .ZN(n1315));
  XNOR2_X1  g0972(.A(n1315), .B(n1314), .ZN(n1316));
  XNOR2_X1  g0973(.A(n1316), .B(n1312), .ZN(n1317));
  XNOR2_X1  g0974(.A(n1317), .B(n1310), .ZN(n1318));
  XNOR2_X1  g0975(.A(n1318), .B(n329), .ZN(n1319));
  XNOR2_X1  g0976(.A(n1319), .B(n453), .ZN(n1320));
  XNOR2_X1  g0977(.A(n1320), .B(n460), .ZN(n1321));
  XNOR2_X1  g0978(.A(n1321), .B(n456), .ZN(n1322));
  XNOR2_X1  g0979(.A(n1322), .B(n467), .ZN(n1323));
  AOI22_X1  g0980(.A1(n1308), .A2(n1307), .B1(367), .B2(n1323), .ZN(n1324));
  XOR2_X1   g0981(.A(n826), .B(n822), .ZN(n1325));
  XNOR2_X1  g0982(.A(n1325), .B(n814), .ZN(n1326));
  XNOR2_X1  g0983(.A(n1326), .B(n449), .ZN(n1327));
  XNOR2_X1  g0984(.A(n1327), .B(n443), .ZN(n1328));
  XNOR2_X1  g0985(.A(n1328), .B(n430), .ZN(n1329));
  XNOR2_X1  g0986(.A(n1329), .B(n433), .ZN(n1330));
  NOR3_X1   g0987(.A1(n1330), .A2(n475), .A3(367), .ZN(n1331));
  INV_X1    g0988(.A(n475), .ZN(n1332));
  OAI21_X1  g0989(.A(367), .B1(n526), .B2(n1332), .ZN(n1333));
  NOR2_X1   g0990(.A1(n1333), .A2(n1330), .ZN(n1334));
  XNOR2_X1  g0991(.A(n819), .B(n441), .ZN(n1335));
  XNOR2_X1  g0992(.A(n1335), .B(n810), .ZN(n1336));
  XNOR2_X1  g0993(.A(n1336), .B(n449), .ZN(n1337));
  XNOR2_X1  g0994(.A(n1337), .B(n443), .ZN(n1338));
  XNOR2_X1  g0995(.A(n1338), .B(n430), .ZN(n1339));
  XNOR2_X1  g0996(.A(n1339), .B(n433), .ZN(n1340));
  AOI211_X1 g0997(.A(n1332), .B(n1340), .C1(n526), .C2(367), .ZN(n1341));
  NOR3_X1   g0998(.A1(n1341), .A2(n1334), .A3(n1331), .ZN(n1342));
  XNOR2_X1  g0999(.A(n1342), .B(n1324), .ZN(11342));
  BUF_X1    g1000(.A(\1 ), .ZN(387));
  BUF_X1    g1001(.A(\1 ), .ZN(388));
  BUF_X1    g1002(.A(248), .ZN(478));
  BUF_X1    g1003(.A(254), .ZN(482));
  BUF_X1    g1004(.A(257), .ZN(484));
  BUF_X1    g1005(.A(260), .ZN(486));
  BUF_X1    g1006(.A(263), .ZN(489));
  BUF_X1    g1007(.A(267), .ZN(492));
  BUF_X1    g1008(.A(274), .ZN(501));
  BUF_X1    g1009(.A(280), .ZN(505));
  BUF_X1    g1010(.A(283), .ZN(507));
  BUF_X1    g1011(.A(286), .ZN(509));
  BUF_X1    g1012(.A(289), .ZN(511));
  BUF_X1    g1013(.A(293), .ZN(513));
  BUF_X1    g1014(.A(296), .ZN(515));
  BUF_X1    g1015(.A(299), .ZN(517));
  BUF_X1    g1016(.A(303), .ZN(519));
  BUF_X1    g1017(.A(307), .ZN(535));
  BUF_X1    g1018(.A(310), .ZN(537));
  BUF_X1    g1019(.A(313), .ZN(539));
  BUF_X1    g1020(.A(316), .ZN(541));
  BUF_X1    g1021(.A(319), .ZN(543));
  BUF_X1    g1022(.A(322), .ZN(545));
  BUF_X1    g1023(.A(325), .ZN(547));
  BUF_X1    g1024(.A(328), .ZN(549));
  BUF_X1    g1025(.A(331), .ZN(551));
  BUF_X1    g1026(.A(334), .ZN(553));
  BUF_X1    g1027(.A(337), .ZN(556));
  BUF_X1    g1028(.A(343), .ZN(559));
  BUF_X1    g1029(.A(346), .ZN(561));
  BUF_X1    g1030(.A(349), .ZN(563));
  BUF_X1    g1031(.A(352), .ZN(565));
  BUF_X1    g1032(.A(355), .ZN(567));
  BUF_X1    g1033(.A(358), .ZN(569));
  BUF_X1    g1034(.A(361), .ZN(571));
  BUF_X1    g1035(.A(364), .ZN(573));
  BUF_X1    g1036(.A(251), .ZN(643));
  BUF_X1    g1037(.A(277), .ZN(707));
  BUF_X1    g1038(.A(340), .ZN(813));
  BUF_X1    g1039(.A(\1 ), .ZN(889));
  BUF_X1    g1040(.A(106), .ZN(945));
  INV_X1    g1041(.A(15), .ZN(1111));
  NAND2_X1  g1042(.A1(242), .A2(n321), .ZN(1112));
  INV_X1    g1043(.A(15), .ZN(1114));
  NAND3_X1  g1044(.A1(134), .A2(133), .A3(n321), .ZN(1489));
  BUF_X1    g1045(.A(\1 ), .ZN(1490));
  NAND3_X1  g1046(.A1(n764), .A2(n720), .A3(n629), .ZN(10103));
  MUX2_X1   g1047(.S(n1053), .B(n1131), .A(n1129), .ZN(10838));
  XNOR2_X1  g1048(.A(n1053), .B(n335), .ZN(10840));
endmodule


