// Benchmark "c880" written by ABC on Wed Oct 05 14:29:36 2022

module c880 ( 
    \1 , 8, 13, 17, 26, 29, 36, 42, 51, 55, 59, 68, 72, 73, 74, 75, 80, 85,
    86, 87, 88, 89, 90, 91, 96, 101, 106, 111, 116, 121, 126, 130, 135,
    138, 143, 146, 149, 152, 153, 156, 159, 165, 171, 177, 183, 189, 195,
    201, 207, 210, 219, 228, 237, 246, 255, 259, 260, 261, 267, 268,
    388, 389, 390, 391, 418, 419, 420, 421, 422, 423, 446, 447, 448, 449,
    450, 767, 768, 850, 863, 864, 865, 866, 874, 878, 879, 880  );
  input  \1 , 8, 13, 17, 26, 29, 36, 42, 51, 55, 59, 68, 72, 73, 74, 75,
    80, 85, 86, 87, 88, 89, 90, 91, 96, 101, 106, 111, 116, 121, 126, 130,
    135, 138, 143, 146, 149, 152, 153, 156, 159, 165, 171, 177, 183, 189,
    195, 201, 207, 210, 219, 228, 237, 246, 255, 259, 260, 261, 267, 268;
  output 388, 389, 390, 391, 418, 419, 420, 421, 422, 423, 446, 447, 448, 449,
    450, 767, 768, 850, 863, 864, 865, 866, 874, 878, 879, 880;
  wire n91, n92, n97, n101, n105, n106, n107, n108, n109, n110, n111, n112,
    n114, n115, n116, n117, n118, n119, n120, n121, n123, n124, n125, n126,
    n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
    n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
    n151, n152, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
    n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
    n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
    n188, n189, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
    n201, n203, n204, n205, n206, n207, n208, n209, n210, n212, n213, n214,
    n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
    n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
    n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n250, n251,
    n252, n253, n254, n255, n256, n257, n258, n259, n261, n262, n263, n264,
    n265, n266, n267, n269, n270, n271, n272, n273, n274, n275, n276, n277,
    n278, n279, n280, n282, n283, n284, n285, n286, n287, n288, n289, n290;
  AND3_X1   g000(.A1(75), .A2(42), .A3(29), .ZN(388));
  AND3_X1   g001(.A1(80), .A2(36), .A3(29), .ZN(389));
  AND3_X1   g002(.A1(42), .A2(36), .A3(29), .ZN(390));
  AND2_X1   g003(.A1(86), .A2(85), .ZN(391));
  AND4_X1   g004(.A1(13), .A2(8), .A3(\1 ), .A4(17), .ZN(418));
  AND4_X1   g005(.A1(17), .A2(13), .A3(\1 ), .A4(26), .ZN(n91));
  INV_X1    g006(.A(n91), .ZN(n92));
  OR2_X1    g007(.A1(n92), .A2(390), .ZN(419));
  NAND3_X1  g008(.A1(80), .A2(75), .A3(59), .ZN(420));
  NAND3_X1  g009(.A1(80), .A2(59), .A3(36), .ZN(421));
  NAND3_X1  g010(.A1(59), .A2(42), .A3(36), .ZN(422));
  OR2_X1    g011(.A1(88), .A2(87), .ZN(n97));
  AND2_X1   g012(.A1(n97), .A2(90), .ZN(423));
  NAND2_X1  g013(.A1(n91), .A2(390), .ZN(446));
  AND3_X1   g014(.A1(51), .A2(26), .A3(\1 ), .ZN(447));
  AND4_X1   g015(.A1(13), .A2(8), .A3(\1 ), .A4(55), .ZN(n101));
  AND3_X1   g016(.A1(n101), .A2(68), .A3(29), .ZN(448));
  AND4_X1   g017(.A1(74), .A2(68), .A3(59), .A4(n101), .ZN(449));
  AND2_X1   g018(.A1(n97), .A2(89), .ZN(450));
  XNOR2_X1  g019(.A(96), .B(91), .ZN(n105));
  XOR2_X1   g020(.A(106), .B(101), .ZN(n106));
  XNOR2_X1  g021(.A(n106), .B(n105), .ZN(n107));
  XNOR2_X1  g022(.A(n107), .B(130), .ZN(n108));
  XNOR2_X1  g023(.A(116), .B(111), .ZN(n109));
  XOR2_X1   g024(.A(126), .B(121), .ZN(n110));
  XOR2_X1   g025(.A(n110), .B(n109), .ZN(n111));
  XNOR2_X1  g026(.A(n111), .B(135), .ZN(n112));
  XNOR2_X1  g027(.A(n112), .B(n108), .ZN(767));
  XNOR2_X1  g028(.A(165), .B(159), .ZN(n114));
  XOR2_X1   g029(.A(177), .B(171), .ZN(n115));
  XNOR2_X1  g030(.A(n115), .B(n114), .ZN(n116));
  XNOR2_X1  g031(.A(n116), .B(130), .ZN(n117));
  XNOR2_X1  g032(.A(189), .B(183), .ZN(n118));
  XOR2_X1   g033(.A(201), .B(195), .ZN(n119));
  XOR2_X1   g034(.A(n119), .B(n118), .ZN(n120));
  XNOR2_X1  g035(.A(n120), .B(207), .ZN(n121));
  XNOR2_X1  g036(.A(n121), .B(n117), .ZN(768));
  INV_X1    g037(.A(153), .ZN(n123));
  INV_X1    g038(.A(17), .ZN(n124));
  NAND3_X1  g039(.A1(51), .A2(26), .A3(\1 ), .ZN(n125));
  AND2_X1   g040(.A1(156), .A2(59), .ZN(n126));
  OR3_X1    g041(.A1(n126), .A2(n125), .A3(n124), .ZN(n127));
  AOI21_X1  g042(.A(n123), .B1(n127), .B2(\1 ), .ZN(n128));
  INV_X1    g043(.A(268), .ZN(n129));
  AND3_X1   g044(.A1(80), .A2(75), .A3(29), .ZN(n130));
  AND4_X1   g045(.A1(447), .A2(n129), .A3(55), .A4(n130), .ZN(n131));
  INV_X1    g046(.A(126), .ZN(n132));
  OR2_X1    g047(.A1(42), .A2(17), .ZN(n133));
  NAND2_X1  g048(.A1(42), .A2(17), .ZN(n134));
  NAND4_X1  g049(.A1(n133), .A2(n126), .A3(447), .A4(n134), .ZN(n135));
  AND3_X1   g050(.A1(75), .A2(59), .A3(42), .ZN(n136));
  NAND4_X1  g051(.A1(17), .A2(8), .A3(\1 ), .A4(51), .ZN(n137));
  OR2_X1    g052(.A1(n137), .A2(n136), .ZN(n138));
  AOI21_X1  g053(.A(n132), .B1(n138), .B2(n135), .ZN(n139));
  NOR3_X1   g054(.A1(n139), .A2(n131), .A3(n128), .ZN(n140));
  XNOR2_X1  g055(.A(n140), .B(201), .ZN(n141));
  NOR2_X1   g056(.A1(n141), .A2(261), .ZN(n142));
  NAND2_X1  g057(.A1(n141), .A2(261), .ZN(n143));
  NAND2_X1  g058(.A1(n143), .A2(219), .ZN(n144));
  INV_X1    g059(.A(201), .ZN(n145));
  NOR2_X1   g060(.A1(n140), .A2(n145), .ZN(n146));
  INV_X1    g061(.A(246), .ZN(n147));
  AND3_X1   g062(.A1(72), .A2(68), .A3(42), .ZN(n148));
  NAND4_X1  g063(.A1(n101), .A2(73), .A3(59), .A4(n148), .ZN(n149));
  AOI22_X1  g064(.A1(255), .A2(267), .B1(210), .B2(121), .ZN(n150));
  OAI221_X1 g065(.A(n150), .B1(n140), .B2(n147), .C1(n145), .C2(n149), .ZN(n151));
  AOI221_X1 g066(.A(n151), .B1(n146), .B2(237), .C1(228), .C2(n141), .ZN(n152));
  OAI21_X1  g067(.A(n152), .B1(n144), .B2(n142), .ZN(850));
  NAND2_X1  g068(.A1(n138), .A2(n135), .ZN(n154));
  INV_X1    g069(.A(143), .ZN(n155));
  AOI21_X1  g070(.A(n155), .B1(n127), .B2(\1 ), .ZN(n156));
  AOI211_X1 g071(.A(n131), .B(n156), .C1(n154), .C2(111), .ZN(n157));
  XNOR2_X1  g072(.A(n157), .B(183), .ZN(n158));
  INV_X1    g073(.A(146), .ZN(n159));
  AOI21_X1  g074(.A(n159), .B1(n127), .B2(\1 ), .ZN(n160));
  INV_X1    g075(.A(116), .ZN(n161));
  AOI21_X1  g076(.A(n161), .B1(n138), .B2(n135), .ZN(n162));
  NOR4_X1   g077(.A1(n160), .A2(n131), .A3(189), .A4(n162), .ZN(n163));
  INV_X1    g078(.A(149), .ZN(n164));
  AOI21_X1  g079(.A(n164), .B1(n127), .B2(\1 ), .ZN(n165));
  INV_X1    g080(.A(121), .ZN(n166));
  AOI21_X1  g081(.A(n166), .B1(n138), .B2(n135), .ZN(n167));
  NOR4_X1   g082(.A1(n165), .A2(n131), .A3(195), .A4(n167), .ZN(n168));
  NOR4_X1   g083(.A1(n163), .A2(n140), .A3(n145), .A4(n168), .ZN(n169));
  INV_X1    g084(.A(261), .ZN(n170));
  NOR4_X1   g085(.A1(n131), .A2(n128), .A3(201), .A4(n139), .ZN(n171));
  NOR4_X1   g086(.A1(n163), .A2(n171), .A3(n170), .A4(n168), .ZN(n172));
  INV_X1    g087(.A(189), .ZN(n173));
  NOR3_X1   g088(.A1(n162), .A2(n160), .A3(n131), .ZN(n174));
  NOR2_X1   g089(.A1(n174), .A2(n173), .ZN(n175));
  INV_X1    g090(.A(195), .ZN(n176));
  NOR3_X1   g091(.A1(n167), .A2(n165), .A3(n131), .ZN(n177));
  NOR3_X1   g092(.A1(n177), .A2(n163), .A3(n176), .ZN(n178));
  OR4_X1    g093(.A1(n175), .A2(n172), .A3(n169), .A4(n178), .ZN(n179));
  NOR2_X1   g094(.A1(n179), .A2(n158), .ZN(n180));
  INV_X1    g095(.A(n158), .ZN(n181));
  NOR4_X1   g096(.A1(n175), .A2(n172), .A3(n169), .A4(n178), .ZN(n182));
  OAI21_X1  g097(.A(219), .B1(n182), .B2(n181), .ZN(n183));
  INV_X1    g098(.A(183), .ZN(n184));
  OR2_X1    g099(.A1(n157), .A2(n184), .ZN(n185));
  INV_X1    g100(.A(n185), .ZN(n186));
  NAND2_X1  g101(.A1(210), .A2(106), .ZN(n187));
  OAI221_X1 g102(.A(n187), .B1(n149), .B2(n184), .C1(n147), .C2(n157), .ZN(n188));
  AOI221_X1 g103(.A(n188), .B1(n186), .B2(237), .C1(228), .C2(n158), .ZN(n189));
  OAI21_X1  g104(.A(n189), .B1(n183), .B2(n180), .ZN(863));
  NOR2_X1   g105(.A1(n177), .A2(n176), .ZN(n191));
  XNOR2_X1  g106(.A(n174), .B(189), .ZN(n192));
  NOR3_X1   g107(.A1(n168), .A2(n171), .A3(n170), .ZN(n193));
  NOR3_X1   g108(.A1(n168), .A2(n140), .A3(n145), .ZN(n194));
  NOR4_X1   g109(.A1(n193), .A2(n192), .A3(n191), .A4(n194), .ZN(n195));
  INV_X1    g110(.A(n192), .ZN(n196));
  NOR3_X1   g111(.A1(n194), .A2(n193), .A3(n191), .ZN(n197));
  OAI21_X1  g112(.A(219), .B1(n197), .B2(n196), .ZN(n198));
  AOI22_X1  g113(.A1(255), .A2(259), .B1(210), .B2(111), .ZN(n199));
  OAI221_X1 g114(.A(n199), .B1(n149), .B2(n173), .C1(n147), .C2(n174), .ZN(n200));
  AOI221_X1 g115(.A(n200), .B1(n175), .B2(237), .C1(228), .C2(n192), .ZN(n201));
  OAI21_X1  g116(.A(n201), .B1(n198), .B2(n195), .ZN(864));
  NOR2_X1   g117(.A1(n171), .A2(n170), .ZN(n203));
  XNOR2_X1  g118(.A(n177), .B(195), .ZN(n204));
  NOR3_X1   g119(.A1(n204), .A2(n203), .A3(n146), .ZN(n205));
  OAI21_X1  g120(.A(n204), .B1(n203), .B2(n146), .ZN(n206));
  NAND2_X1  g121(.A1(n206), .A2(219), .ZN(n207));
  AOI22_X1  g122(.A1(255), .A2(260), .B1(210), .B2(116), .ZN(n208));
  OAI221_X1 g123(.A(n208), .B1(n149), .B2(n176), .C1(n147), .C2(n177), .ZN(n209));
  AOI221_X1 g124(.A(n209), .B1(n191), .B2(237), .C1(228), .C2(n204), .ZN(n210));
  OAI21_X1  g125(.A(n210), .B1(n207), .B2(n205), .ZN(865));
  INV_X1    g126(.A(159), .ZN(n212));
  INV_X1    g127(.A(91), .ZN(n213));
  AOI21_X1  g128(.A(n213), .B1(n138), .B2(n135), .ZN(n214));
  INV_X1    g129(.A(55), .ZN(n215));
  OR3_X1    g130(.A1(n126), .A2(n125), .A3(n215), .ZN(n216));
  NAND2_X1  g131(.A1(138), .A2(8), .ZN(n217));
  NAND4_X1  g132(.A1(447), .A2(n129), .A3(17), .A4(n130), .ZN(n218));
  OAI211_X1 g133(.A(n217), .B(n218), .C1(n216), .C2(n155), .ZN(n219));
  NOR2_X1   g134(.A1(n219), .A2(n214), .ZN(n220));
  NOR2_X1   g135(.A1(n220), .A2(n212), .ZN(n221));
  INV_X1    g136(.A(n221), .ZN(n222));
  AND2_X1   g137(.A1(n157), .A2(n184), .ZN(n223));
  OAI21_X1  g138(.A(n185), .B1(n182), .B2(n223), .ZN(n224));
  INV_X1    g139(.A(96), .ZN(n225));
  AOI21_X1  g140(.A(n225), .B1(n138), .B2(n135), .ZN(n226));
  NAND2_X1  g141(.A1(138), .A2(51), .ZN(n227));
  OAI211_X1 g142(.A(n218), .B(n227), .C1(n216), .C2(n159), .ZN(n228));
  NOR3_X1   g143(.A1(n228), .A2(n226), .A3(165), .ZN(n229));
  INV_X1    g144(.A(101), .ZN(n230));
  AOI21_X1  g145(.A(n230), .B1(n138), .B2(n135), .ZN(n231));
  NAND2_X1  g146(.A1(138), .A2(17), .ZN(n232));
  OAI211_X1 g147(.A(n218), .B(n232), .C1(n216), .C2(n164), .ZN(n233));
  NOR3_X1   g148(.A1(n233), .A2(n231), .A3(171), .ZN(n234));
  INV_X1    g149(.A(106), .ZN(n235));
  AOI21_X1  g150(.A(n235), .B1(n138), .B2(n135), .ZN(n236));
  NAND2_X1  g151(.A1(152), .A2(138), .ZN(n237));
  OAI211_X1 g152(.A(n218), .B(n237), .C1(n216), .C2(n123), .ZN(n238));
  NOR3_X1   g153(.A1(n238), .A2(n236), .A3(177), .ZN(n239));
  NOR3_X1   g154(.A1(n239), .A2(n234), .A3(n229), .ZN(n240));
  INV_X1    g155(.A(177), .ZN(n241));
  NOR2_X1   g156(.A1(n238), .A2(n236), .ZN(n242));
  NOR4_X1   g157(.A1(n234), .A2(n229), .A3(n241), .A4(n242), .ZN(n243));
  OAI21_X1  g158(.A(165), .B1(n228), .B2(n226), .ZN(n244));
  OAI21_X1  g159(.A(171), .B1(n233), .B2(n231), .ZN(n245));
  OAI21_X1  g160(.A(n244), .B1(n245), .B2(n229), .ZN(n246));
  AOI211_X1 g161(.A(n243), .B(n246), .C1(n240), .C2(n224), .ZN(n247));
  NOR3_X1   g162(.A1(n219), .A2(n214), .A3(159), .ZN(n248));
  OAI21_X1  g163(.A(n222), .B1(n248), .B2(n247), .ZN(866));
  INV_X1    g164(.A(228), .ZN(n250));
  XNOR2_X1  g165(.A(n242), .B(n241), .ZN(n251));
  INV_X1    g166(.A(n223), .ZN(n252));
  AOI21_X1  g167(.A(n186), .B1(n179), .B2(n252), .ZN(n253));
  AND2_X1   g168(.A1(n251), .A2(n253), .ZN(n254));
  OAI21_X1  g169(.A(219), .B1(n251), .B2(n253), .ZN(n255));
  NOR2_X1   g170(.A1(n242), .A2(n241), .ZN(n256));
  NAND2_X1  g171(.A1(210), .A2(101), .ZN(n257));
  OAI221_X1 g172(.A(n257), .B1(n149), .B2(n241), .C1(n147), .C2(n242), .ZN(n258));
  AOI21_X1  g173(.A(n258), .B1(n256), .B2(237), .ZN(n259));
  OAI221_X1 g174(.A(n259), .B1(n254), .B2(n255), .C1(n251), .C2(n250), .ZN(874));
  XNOR2_X1  g175(.A(n220), .B(n212), .ZN(n261));
  AND2_X1   g176(.A1(n261), .A2(n247), .ZN(n262));
  OAI21_X1  g177(.A(219), .B1(n261), .B2(n247), .ZN(n263));
  INV_X1    g178(.A(210), .ZN(n264));
  OAI21_X1  g179(.A(246), .B1(n219), .B2(n214), .ZN(n265));
  OAI221_X1 g180(.A(n265), .B1(n129), .B2(n264), .C1(n212), .C2(n149), .ZN(n266));
  AOI21_X1  g181(.A(n266), .B1(n221), .B2(237), .ZN(n267));
  OAI221_X1 g182(.A(n267), .B1(n262), .B2(n263), .C1(n261), .C2(n250), .ZN(878));
  INV_X1    g183(.A(n244), .ZN(n269));
  OR2_X1    g184(.A1(n269), .A2(n229), .ZN(n270));
  INV_X1    g185(.A(n245), .ZN(n271));
  NOR2_X1   g186(.A1(n239), .A2(n234), .ZN(n272));
  NOR3_X1   g187(.A1(n242), .A2(n234), .A3(n241), .ZN(n273));
  AOI211_X1 g188(.A(n271), .B(n273), .C1(n272), .C2(n224), .ZN(n274));
  AND2_X1   g189(.A1(n274), .A2(n270), .ZN(n275));
  OAI21_X1  g190(.A(219), .B1(n274), .B2(n270), .ZN(n276));
  INV_X1    g191(.A(165), .ZN(n277));
  OAI21_X1  g192(.A(246), .B1(n228), .B2(n226), .ZN(n278));
  OAI221_X1 g193(.A(n278), .B1(n264), .B2(n213), .C1(n277), .C2(n149), .ZN(n279));
  AOI21_X1  g194(.A(n279), .B1(n269), .B2(237), .ZN(n280));
  OAI221_X1 g195(.A(n280), .B1(n275), .B2(n276), .C1(n270), .C2(n250), .ZN(879));
  OR2_X1    g196(.A1(n233), .A2(n231), .ZN(n282));
  XNOR2_X1  g197(.A(n282), .B(171), .ZN(n283));
  INV_X1    g198(.A(n239), .ZN(n284));
  AOI21_X1  g199(.A(n256), .B1(n284), .B2(n224), .ZN(n285));
  AND2_X1   g200(.A1(n285), .A2(n283), .ZN(n286));
  OAI21_X1  g201(.A(219), .B1(n285), .B2(n283), .ZN(n287));
  INV_X1    g202(.A(171), .ZN(n288));
  OAI22_X1  g203(.A1(n264), .A2(n225), .B1(n288), .B2(n149), .ZN(n289));
  AOI221_X1 g204(.A(n289), .B1(n282), .B2(246), .C1(237), .C2(n271), .ZN(n290));
  OAI221_X1 g205(.A(n290), .B1(n286), .B2(n287), .C1(n283), .C2(n250), .ZN(880));
endmodule


