// Benchmark "c432" written by ABC on Tue Nov 29 09:37:14 2022

module c432 ( 
    1, 4, 8, 11, 14, 17, 21, 24, 27, 30, 34, 37, 40, 43, 47, 50, 53, 56,
    60, 63, 66, 69, 73, 76, 79, 82, 86, 89, 92, 95, 99, 102, 105, 108, 112,
    115,
    223, 329, 370, 421, 430, 431, 432  );
  input  1, 4, 8, 11, 14, 17, 21, 24, 27, 30, 34, 37, 40, 43, 47, 50,
    53, 56, 60, 63, 66, 69, 73, 76, 79, 82, 86, 89, 92, 95, 99, 102, 105,
    108, 112, 115;
  output 223, 329, 370, 421, 430, 431, 432;
  wire n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
    n57, n58, n59, n60, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
    n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n88,
    n89, n90, n94, n95, n96, n97, n99, n100, n101, n102, n103, n105, n106,
    n107, n108, n111, n116, n117, n118, n119, n120, n121, n122, n123, n124,
    n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
    n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
    n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
    n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
    n174, n175, n177, n178, n179, n180, n181, n182, n183, n184, n186, n187,
    n189, n190, n191;
  INV_X1    g000(.A(108), .ZN(n43));
  NOR2_X1   g001(.A1(n43), .A2(102), .ZN(n44));
  INV_X1    g002(.A(82), .ZN(n45));
  INV_X1    g003(.A(95), .ZN(n46));
  OAI22_X1  g004(.A1(89), .A2(n46), .B1(n45), .B2(76), .ZN(n47));
  NOR2_X1   g005(.A1(n47), .A2(n44), .ZN(n48));
  INV_X1    g006(.A(4), .ZN(n49));
  INV_X1    g007(.A(17), .ZN(n50));
  OAI22_X1  g008(.A1(11), .A2(n50), .B1(n49), .B2(1), .ZN(n51));
  INV_X1    g009(.A(43), .ZN(n52));
  NOR2_X1   g010(.A1(n52), .A2(37), .ZN(n53));
  INV_X1    g011(.A(30), .ZN(n54));
  NOR2_X1   g012(.A1(n54), .A2(24), .ZN(n55));
  INV_X1    g013(.A(56), .ZN(n56));
  INV_X1    g014(.A(69), .ZN(n57));
  OAI22_X1  g015(.A1(63), .A2(n57), .B1(n56), .B2(50), .ZN(n58));
  NOR4_X1   g016(.A1(n55), .A2(n53), .A3(n51), .A4(n58), .ZN(n59));
  AND2_X1   g017(.A1(n59), .A2(n48), .ZN(n60));
  INV_X1    g018(.A(n60), .ZN(223));
  INV_X1    g019(.A(112), .ZN(n62));
  OR4_X1    g020(.A1(n55), .A2(n53), .A3(n51), .A4(n58), .ZN(n63));
  OAI22_X1  g021(.A1(n47), .A2(n63), .B1(n43), .B2(102), .ZN(n64));
  NAND3_X1  g022(.A1(n64), .A2(n62), .A3(108), .ZN(n65));
  NOR2_X1   g023(.A1(n46), .A2(89), .ZN(n66));
  XNOR2_X1  g024(.A(n60), .B(n66), .ZN(n67));
  NOR2_X1   g025(.A1(99), .A2(n46), .ZN(n68));
  INV_X1    g026(.A(n68), .ZN(n69));
  NOR2_X1   g027(.A1(n45), .A2(76), .ZN(n70));
  XNOR2_X1  g028(.A(n60), .B(n70), .ZN(n71));
  NOR2_X1   g029(.A1(86), .A2(n45), .ZN(n72));
  INV_X1    g030(.A(n72), .ZN(n73));
  OAI221_X1 g031(.A(n65), .B1(n69), .B2(n67), .C1(n73), .C2(n71), .ZN(n74));
  NOR2_X1   g032(.A1(n49), .A2(1), .ZN(n75));
  XOR2_X1   g033(.A(n60), .B(n75), .Z(n76));
  NOR2_X1   g034(.A1(8), .A2(n49), .ZN(n77));
  AND2_X1   g035(.A1(n77), .A2(n76), .ZN(n78));
  NOR2_X1   g036(.A1(n50), .A2(11), .ZN(n79));
  XOR2_X1   g037(.A(n60), .B(n79), .Z(n80));
  NOR2_X1   g038(.A1(21), .A2(n50), .ZN(n81));
  AND2_X1   g039(.A1(n81), .A2(n80), .ZN(n82));
  INV_X1    g040(.A(47), .ZN(n83));
  INV_X1    g041(.A(37), .ZN(n84));
  OAI211_X1 g042(.A(n83), .B(43), .C1(n60), .C2(n53), .ZN(n88));
  INV_X1    g043(.A(34), .ZN(n89));
  INV_X1    g044(.A(24), .ZN(n90));
  OAI211_X1 g045(.A(n89), .B(30), .C1(n60), .C2(n55), .ZN(n94));
  INV_X1    g046(.A(73), .ZN(n95));
  INV_X1    g047(.A(63), .ZN(n96));
  NAND2_X1  g048(.A1(69), .A2(n96), .ZN(n97));
  AOI21_X1  g049(.A(n97), .B1(n59), .B2(n48), .ZN(n99));
  OAI211_X1 g050(.A(n95), .B(69), .C1(n60), .C2(n99), .ZN(n100));
  INV_X1    g051(.A(60), .ZN(n101));
  INV_X1    g052(.A(50), .ZN(n102));
  NAND2_X1  g053(.A1(56), .A2(n102), .ZN(n103));
  AOI21_X1  g054(.A(n103), .B1(n59), .B2(n48), .ZN(n105));
  OAI211_X1 g055(.A(n101), .B(56), .C1(n60), .C2(n105), .ZN(n106));
  NAND4_X1  g056(.A1(n100), .A2(n94), .A3(n88), .A4(n106), .ZN(n107));
  NOR4_X1   g057(.A1(n82), .A2(n78), .A3(n74), .A4(n107), .ZN(n108));
  INV_X1    g058(.A(n108), .ZN(329));
  XOR2_X1   g059(.A(n60), .B(n70), .Z(n111));
  NOR2_X1   g060(.A1(112), .A2(n43), .ZN(n116));
  AND2_X1   g061(.A1(n116), .A2(n64), .ZN(n117));
  NOR2_X1   g062(.A1(115), .A2(n43), .ZN(n118));
  OAI211_X1 g063(.A(n64), .B(n118), .C1(n117), .C2(n108), .ZN(n119));
  NOR2_X1   g064(.A1(n69), .A2(n67), .ZN(n120));
  XNOR2_X1  g065(.A(n108), .B(n120), .ZN(n121));
  OR3_X1    g066(.A1(n67), .A2(105), .A3(n46), .ZN(n122));
  NOR2_X1   g067(.A1(n73), .A2(n71), .ZN(n123));
  XNOR2_X1  g068(.A(n108), .B(n123), .ZN(n124));
  INV_X1    g069(.A(92), .ZN(n125));
  NAND3_X1  g070(.A1(n111), .A2(n125), .A3(82), .ZN(n126));
  OAI221_X1 g071(.A(n119), .B1(n122), .B2(n121), .C1(n126), .C2(n124), .ZN(n127));
  XNOR2_X1  g072(.A(n108), .B(n78), .ZN(n128));
  NOR2_X1   g073(.A1(14), .A2(n49), .ZN(n129));
  NAND2_X1  g074(.A1(n129), .A2(n76), .ZN(n130));
  XNOR2_X1  g075(.A(n108), .B(n82), .ZN(n131));
  INV_X1    g076(.A(27), .ZN(n132));
  NAND3_X1  g077(.A1(n80), .A2(n132), .A3(17), .ZN(n133));
  OAI22_X1  g078(.A1(n131), .A2(n133), .B1(n130), .B2(n128), .ZN(n134));
  XOR2_X1   g079(.A(n108), .B(n88), .Z(n135));
  INV_X1    g080(.A(53), .ZN(n136));
  OAI211_X1 g081(.A(n136), .B(43), .C1(n60), .C2(n53), .ZN(n137));
  XOR2_X1   g082(.A(n108), .B(n94), .Z(n138));
  INV_X1    g083(.A(40), .ZN(n139));
  OAI211_X1 g084(.A(n139), .B(30), .C1(n60), .C2(n55), .ZN(n140));
  OAI22_X1  g085(.A1(n138), .A2(n140), .B1(n137), .B2(n135), .ZN(n141));
  XOR2_X1   g086(.A(n108), .B(n100), .Z(n142));
  NOR2_X1   g087(.A1(79), .A2(n57), .ZN(n143));
  OAI21_X1  g088(.A(n143), .B1(n99), .B2(n60), .ZN(n144));
  XOR2_X1   g089(.A(n108), .B(n106), .Z(n145));
  INV_X1    g090(.A(66), .ZN(n146));
  OAI211_X1 g091(.A(n146), .B(56), .C1(n60), .C2(n105), .ZN(n147));
  OAI22_X1  g092(.A1(n145), .A2(n147), .B1(n144), .B2(n142), .ZN(n148));
  OR4_X1    g093(.A1(n141), .A2(n134), .A3(n127), .A4(n148), .ZN(370));
  NAND2_X1  g094(.A1(370), .A2(14), .ZN(n150));
  AOI221_X1 g095(.A(n49), .B1(8), .B2(329), .C1(1), .C2(223), .ZN(n151));
  OAI221_X1 g096(.A(56), .B1(n101), .B2(n108), .C1(n102), .C2(n60), .ZN(n152));
  AOI21_X1  g097(.A(n152), .B1(370), .B2(66), .ZN(n153));
  OAI221_X1 g098(.A(43), .B1(n83), .B2(n108), .C1(n84), .C2(n60), .ZN(n154));
  AOI21_X1  g099(.A(n154), .B1(370), .B2(53), .ZN(n155));
  INV_X1    g100(.A(86), .ZN(n156));
  AOI21_X1  g101(.A(n45), .B1(223), .B2(76), .ZN(n157));
  OAI21_X1  g102(.A(n157), .B1(n108), .B2(n156), .ZN(n158));
  AOI21_X1  g103(.A(n158), .B1(370), .B2(92), .ZN(n159));
  OAI221_X1 g104(.A(69), .B1(n95), .B2(n108), .C1(n96), .C2(n60), .ZN(n160));
  AOI21_X1  g105(.A(n160), .B1(370), .B2(79), .ZN(n161));
  NOR4_X1   g106(.A1(n159), .A2(n155), .A3(n153), .A4(n161), .ZN(n162));
  INV_X1    g107(.A(21), .ZN(n163));
  AOI21_X1  g108(.A(n50), .B1(223), .B2(11), .ZN(n164));
  OAI21_X1  g109(.A(n164), .B1(n108), .B2(n163), .ZN(n165));
  AOI21_X1  g110(.A(n165), .B1(370), .B2(27), .ZN(n166));
  OAI221_X1 g111(.A(30), .B1(n89), .B2(n108), .C1(n90), .C2(n60), .ZN(n167));
  AOI21_X1  g112(.A(n167), .B1(370), .B2(40), .ZN(n168));
  AOI21_X1  g113(.A(n43), .B1(223), .B2(102), .ZN(n169));
  OAI21_X1  g114(.A(n169), .B1(n108), .B2(n62), .ZN(n170));
  AOI21_X1  g115(.A(n170), .B1(370), .B2(115), .ZN(n171));
  INV_X1    g116(.A(89), .ZN(n172));
  OAI21_X1  g117(.A(95), .B1(n60), .B2(n172), .ZN(n173));
  AOI221_X1 g118(.A(n173), .B1(329), .B2(99), .C1(105), .C2(370), .ZN(n174));
  NOR4_X1   g119(.A1(n171), .A2(n168), .A3(n166), .A4(n174), .ZN(n175));
  AOI22_X1  g120(.A1(n162), .A2(n175), .B1(n151), .B2(n150), .ZN(421));
  NOR4_X1   g121(.A1(n141), .A2(n134), .A3(n127), .A4(n148), .ZN(n177));
  INV_X1    g122(.A(n152), .ZN(n178));
  OAI21_X1  g123(.A(n178), .B1(n177), .B2(n146), .ZN(n179));
  INV_X1    g124(.A(n154), .ZN(n180));
  OAI21_X1  g125(.A(n180), .B1(n177), .B2(n136), .ZN(n181));
  OAI221_X1 g126(.A(n164), .B1(n108), .B2(n163), .C1(n132), .C2(n177), .ZN(n182));
  INV_X1    g127(.A(n167), .ZN(n183));
  OAI21_X1  g128(.A(n183), .B1(n177), .B2(n139), .ZN(n184));
  NAND4_X1  g129(.A1(n182), .A2(n181), .A3(n179), .A4(n184), .ZN(430));
  NAND4_X1  g130(.A1(n161), .A2(n181), .A3(n179), .A4(n184), .ZN(n186));
  NAND3_X1  g131(.A1(n159), .A2(n181), .A3(n179), .ZN(n187));
  NAND4_X1  g132(.A1(n186), .A2(n184), .A3(n182), .A4(n187), .ZN(431));
  OAI221_X1 g133(.A(n157), .B1(n108), .B2(n156), .C1(n125), .C2(n177), .ZN(n189));
  NAND4_X1  g134(.A1(n184), .A2(n189), .A3(n181), .A4(n174), .ZN(n190));
  AOI21_X1  g135(.A(n166), .B1(n184), .B2(n155), .ZN(n191));
  NAND3_X1  g136(.A1(n191), .A2(n190), .A3(n186), .ZN(432));
endmodule


