// Benchmark "c6288" written by ABC on Wed Oct 05 14:34:49 2022

module c6288 ( 
    \1 , 18, 35, 52, 69, 86, 103, 120, 137, 154, 171, 188, 205, 222, 239,
    256, 273, 290, 307, 324, 341, 358, 375, 392, 409, 426, 443, 460, 477,
    494, 511, 528,
    545, 1581, 1901, 2223, 2548, 2877, 3211, 3552, 3895, 4241, 4591, 4946,
    5308, 5672, 5971, 6123, 6150, 6160, 6170, 6180, 6190, 6200, 6210, 6220,
    6230, 6240, 6250, 6260, 6270, 6280, 6287, 6288  );
  input  \1 , 18, 35, 52, 69, 86, 103, 120, 137, 154, 171, 188, 205, 222,
    239, 256, 273, 290, 307, 324, 341, 358, 375, 392, 409, 426, 443, 460,
    477, 494, 511, 528;
  output 545, 1581, 1901, 2223, 2548, 2877, 3211, 3552, 3895, 4241, 4591,
    4946, 5308, 5672, 5971, 6123, 6150, 6160, 6170, 6180, 6190, 6200, 6210,
    6220, 6230, 6240, 6250, 6260, 6270, 6280, 6287, 6288;
  wire n65, n66, n68, n69, n70, n71, n72, n74, n75, n76, n77, n78, n79, n80,
    n81, n82, n83, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
    n96, n97, n98, n99, n100, n101, n102, n103, n105, n106, n107, n108,
    n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
    n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
    n133, n134, n135, n136, n138, n139, n140, n141, n142, n143, n144, n145,
    n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
    n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
    n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
    n182, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
    n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
    n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
    n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
    n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n243,
    n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
    n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
    n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
    n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
    n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
    n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n315, n316,
    n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
    n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
    n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
    n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
    n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
    n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
    n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n400, n401,
    n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
    n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
    n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
    n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
    n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
    n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
    n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
    n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n498,
    n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
    n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
    n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
    n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
    n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
    n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
    n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
    n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
    n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
    n607, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
    n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
    n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
    n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
    n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
    n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
    n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
    n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
    n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
    n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
    n728, n729, n730, n731, n733, n734, n735, n736, n737, n738, n739, n740,
    n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
    n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
    n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
    n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
    n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
    n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
    n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
    n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
    n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
    n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
    n861, n862, n863, n864, n865, n866, n867, n868, n870, n871, n872, n873,
    n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
    n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
    n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
    n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
    n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
    n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
    n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
    n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
    n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
    n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
    n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
    n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
    n1015, n1016, n1017, n1018, n1020, n1021, n1022, n1023, n1024, n1025,
    n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
    n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
    n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
    n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
    n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
    n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
    n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
    n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
    n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
    n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
    n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
    n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
    n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
    n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
    n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
    n1176, n1177, n1178, n1179, n1180, n1181, n1183, n1184, n1185, n1186,
    n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
    n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
    n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
    n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
    n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
    n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
    n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
    n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
    n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
    n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
    n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
    n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
    n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
    n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
    n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
    n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
    n1347, n1348, n1349, n1350, n1351, n1352, n1354, n1355, n1356, n1357,
    n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
    n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
    n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
    n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
    n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407,
    n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417,
    n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427,
    n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437,
    n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447,
    n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457,
    n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467,
    n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477,
    n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487,
    n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497,
    n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507,
    n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517,
    n1518, n1519, n1520, n1521, n1522, n1524, n1525, n1526, n1527, n1528,
    n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538,
    n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548,
    n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558,
    n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568,
    n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578,
    n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588,
    n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598,
    n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608,
    n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618,
    n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628,
    n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638,
    n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648,
    n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658,
    n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668,
    n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678,
    n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688,
    n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699,
    n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709,
    n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719,
    n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729,
    n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739,
    n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749,
    n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759,
    n1760, n1761, n1762, n1764, n1765, n1766, n1767, n1768, n1769, n1770,
    n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780,
    n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790,
    n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800,
    n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810,
    n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820,
    n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830,
    n1831, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841,
    n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851,
    n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861,
    n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871,
    n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881,
    n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891,
    n1892, n1893, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
    n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
    n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
    n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
    n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
    n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1952, n1953,
    n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963,
    n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973,
    n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983,
    n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993,
    n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2002, n2003, n2004,
    n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
    n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
    n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
    n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
    n2045, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055,
    n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065,
    n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075,
    n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2085, n2086,
    n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096,
    n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106,
    n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116,
    n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127,
    n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137,
    n2138, n2139, n2140, n2141, n2142, n2144, n2145, n2146, n2147, n2148,
    n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158,
    n2159, n2160, n2161, n2162, n2163, n2165, n2166, n2167, n2168, n2169,
    n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2179, n2180,
    n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188;
  AND2_X1   g0000(.A1(273), .A2(\1 ), .ZN(545));
  AND4_X1   g0001(.A1(273), .A2(18), .A3(\1 ), .A4(290), .ZN(n65));
  AOI22_X1  g0002(.A1(273), .A2(18), .B1(\1 ), .B2(290), .ZN(n66));
  NOR2_X1   g0003(.A1(n66), .A2(n65), .ZN(1581));
  AND4_X1   g0004(.A1(273), .A2(35), .A3(18), .A4(290), .ZN(n68));
  AOI22_X1  g0005(.A1(273), .A2(35), .B1(18), .B2(290), .ZN(n69));
  NOR2_X1   g0006(.A1(n69), .A2(n68), .ZN(n70));
  XOR2_X1   g0007(.A(n70), .B(n65), .ZN(n71));
  NAND2_X1  g0008(.A1(307), .A2(\1 ), .ZN(n72));
  XNOR2_X1  g0009(.A(n72), .B(n71), .ZN(1901));
  AND4_X1   g0010(.A1(273), .A2(52), .A3(35), .A4(290), .ZN(n74));
  AOI22_X1  g0011(.A1(273), .A2(52), .B1(35), .B2(290), .ZN(n75));
  NOR2_X1   g0012(.A1(n75), .A2(n74), .ZN(n76));
  XNOR2_X1  g0013(.A(n76), .B(n68), .ZN(n77));
  AND2_X1   g0014(.A1(307), .A2(18), .ZN(n78));
  XNOR2_X1  g0015(.A(n78), .B(n77), .ZN(n79));
  NOR2_X1   g0016(.A1(n70), .A2(n65), .ZN(n80));
  AOI21_X1  g0017(.A(n80), .B1(n72), .B2(n71), .ZN(n81));
  XOR2_X1   g0018(.A(n81), .B(n79), .ZN(n82));
  NAND2_X1  g0019(.A1(324), .A2(\1 ), .ZN(n83));
  XNOR2_X1  g0020(.A(n83), .B(n82), .ZN(2223));
  AND4_X1   g0021(.A1(273), .A2(69), .A3(52), .A4(290), .ZN(n85));
  AOI22_X1  g0022(.A1(273), .A2(69), .B1(52), .B2(290), .ZN(n86));
  NOR2_X1   g0023(.A1(n86), .A2(n85), .ZN(n87));
  XNOR2_X1  g0024(.A(n87), .B(n74), .ZN(n88));
  AND2_X1   g0025(.A1(307), .A2(35), .ZN(n89));
  XNOR2_X1  g0026(.A(n89), .B(n88), .ZN(n90));
  NOR2_X1   g0027(.A1(n76), .A2(n68), .ZN(n91));
  OAI21_X1  g0028(.A(n68), .B1(n75), .B2(n74), .ZN(n92));
  OR3_X1    g0029(.A1(n75), .A2(n74), .A3(n68), .ZN(n93));
  AOI21_X1  g0030(.A(n78), .B1(n93), .B2(n92), .ZN(n94));
  NOR2_X1   g0031(.A1(n94), .A2(n91), .ZN(n95));
  XNOR2_X1  g0032(.A(n95), .B(n90), .ZN(n96));
  AND2_X1   g0033(.A1(324), .A2(18), .ZN(n97));
  XNOR2_X1  g0034(.A(n97), .B(n96), .ZN(n98));
  NOR2_X1   g0035(.A1(n81), .A2(n79), .ZN(n99));
  AOI21_X1  g0036(.A(n99), .B1(n83), .B2(n82), .ZN(n100));
  XOR2_X1   g0037(.A(n100), .B(n98), .ZN(n101));
  AND2_X1   g0038(.A1(341), .A2(\1 ), .ZN(n102));
  INV_X1    g0039(.A(n102), .ZN(n103));
  XNOR2_X1  g0040(.A(n103), .B(n101), .ZN(2548));
  AND4_X1   g0041(.A1(273), .A2(86), .A3(69), .A4(290), .ZN(n105));
  AOI22_X1  g0042(.A1(273), .A2(86), .B1(69), .B2(290), .ZN(n106));
  NOR2_X1   g0043(.A1(n106), .A2(n105), .ZN(n107));
  XNOR2_X1  g0044(.A(n107), .B(n85), .ZN(n108));
  AND2_X1   g0045(.A1(307), .A2(52), .ZN(n109));
  XNOR2_X1  g0046(.A(n109), .B(n108), .ZN(n110));
  NOR2_X1   g0047(.A1(n87), .A2(n74), .ZN(n111));
  OAI21_X1  g0048(.A(n74), .B1(n86), .B2(n85), .ZN(n112));
  OR3_X1    g0049(.A1(n86), .A2(n85), .A3(n74), .ZN(n113));
  AOI21_X1  g0050(.A(n89), .B1(n113), .B2(n112), .ZN(n114));
  NOR2_X1   g0051(.A1(n114), .A2(n111), .ZN(n115));
  XNOR2_X1  g0052(.A(n115), .B(n110), .ZN(n116));
  AND2_X1   g0053(.A1(324), .A2(35), .ZN(n117));
  XNOR2_X1  g0054(.A(n117), .B(n116), .ZN(n118));
  NOR2_X1   g0055(.A1(n95), .A2(n90), .ZN(n119));
  OR2_X1    g0056(.A1(n76), .A2(n68), .ZN(n120));
  NAND2_X1  g0057(.A1(307), .A2(35), .ZN(n121));
  AOI21_X1  g0058(.A(n121), .B1(n113), .B2(n112), .ZN(n122));
  AND3_X1   g0059(.A1(n121), .A2(n113), .A3(n112), .ZN(n123));
  OAI221_X1 g0060(.A(n120), .B1(n78), .B2(n77), .C1(n123), .C2(n122), .ZN(n124));
  NAND3_X1  g0061(.A1(n121), .A2(n113), .A3(n112), .ZN(n125));
  OAI221_X1 g0062(.A(n125), .B1(n88), .B2(n114), .C1(n94), .C2(n91), .ZN(n126));
  AOI21_X1  g0063(.A(n97), .B1(n126), .B2(n124), .ZN(n127));
  NOR2_X1   g0064(.A1(n127), .A2(n119), .ZN(n128));
  XNOR2_X1  g0065(.A(n128), .B(n118), .ZN(n129));
  AND2_X1   g0066(.A1(341), .A2(18), .ZN(n130));
  XNOR2_X1  g0067(.A(n130), .B(n129), .ZN(n131));
  NOR2_X1   g0068(.A1(n100), .A2(n98), .ZN(n132));
  AOI21_X1  g0069(.A(n132), .B1(n103), .B2(n101), .ZN(n133));
  XOR2_X1   g0070(.A(n133), .B(n131), .ZN(n134));
  AND2_X1   g0071(.A1(358), .A2(\1 ), .ZN(n135));
  INV_X1    g0072(.A(n135), .ZN(n136));
  XNOR2_X1  g0073(.A(n136), .B(n134), .ZN(2877));
  AND4_X1   g0074(.A1(273), .A2(103), .A3(86), .A4(290), .ZN(n138));
  AOI22_X1  g0075(.A1(273), .A2(103), .B1(86), .B2(290), .ZN(n139));
  NOR2_X1   g0076(.A1(n139), .A2(n138), .ZN(n140));
  XNOR2_X1  g0077(.A(n140), .B(n105), .ZN(n141));
  AND2_X1   g0078(.A1(307), .A2(69), .ZN(n142));
  XNOR2_X1  g0079(.A(n142), .B(n141), .ZN(n143));
  NOR2_X1   g0080(.A1(n107), .A2(n85), .ZN(n144));
  OAI21_X1  g0081(.A(n85), .B1(n106), .B2(n105), .ZN(n145));
  OR3_X1    g0082(.A1(n106), .A2(n105), .A3(n85), .ZN(n146));
  AOI21_X1  g0083(.A(n109), .B1(n146), .B2(n145), .ZN(n147));
  NOR2_X1   g0084(.A1(n147), .A2(n144), .ZN(n148));
  XNOR2_X1  g0085(.A(n148), .B(n143), .ZN(n149));
  AND2_X1   g0086(.A1(324), .A2(52), .ZN(n150));
  XNOR2_X1  g0087(.A(n150), .B(n149), .ZN(n151));
  NOR2_X1   g0088(.A1(n115), .A2(n110), .ZN(n152));
  OR2_X1    g0089(.A1(n87), .A2(n74), .ZN(n153));
  NAND2_X1  g0090(.A1(307), .A2(52), .ZN(n154));
  AOI21_X1  g0091(.A(n154), .B1(n146), .B2(n145), .ZN(n155));
  AND3_X1   g0092(.A1(n154), .A2(n146), .A3(n145), .ZN(n156));
  OAI221_X1 g0093(.A(n153), .B1(n89), .B2(n88), .C1(n156), .C2(n155), .ZN(n157));
  NAND3_X1  g0094(.A1(n154), .A2(n146), .A3(n145), .ZN(n158));
  OAI221_X1 g0095(.A(n158), .B1(n108), .B2(n147), .C1(n114), .C2(n111), .ZN(n159));
  AOI21_X1  g0096(.A(n117), .B1(n159), .B2(n157), .ZN(n160));
  NOR2_X1   g0097(.A1(n160), .A2(n152), .ZN(n161));
  XNOR2_X1  g0098(.A(n161), .B(n151), .ZN(n162));
  AND2_X1   g0099(.A1(341), .A2(35), .ZN(n163));
  XNOR2_X1  g0100(.A(n163), .B(n162), .ZN(n164));
  NOR2_X1   g0101(.A1(n128), .A2(n118), .ZN(n165));
  OAI22_X1  g0102(.A1(n122), .A2(n123), .B1(n94), .B2(n91), .ZN(n166));
  INV_X1    g0103(.A(n117), .ZN(n167));
  AOI21_X1  g0104(.A(n167), .B1(n159), .B2(n157), .ZN(n168));
  AND3_X1   g0105(.A1(n167), .A2(n159), .A3(n157), .ZN(n169));
  OAI221_X1 g0106(.A(n166), .B1(n97), .B2(n96), .C1(n169), .C2(n168), .ZN(n170));
  NAND3_X1  g0107(.A1(n167), .A2(n159), .A3(n157), .ZN(n171));
  OAI221_X1 g0108(.A(n171), .B1(n116), .B2(n160), .C1(n127), .C2(n119), .ZN(n172));
  AOI21_X1  g0109(.A(n130), .B1(n172), .B2(n170), .ZN(n173));
  NOR2_X1   g0110(.A1(n173), .A2(n165), .ZN(n174));
  XNOR2_X1  g0111(.A(n174), .B(n164), .ZN(n175));
  AND2_X1   g0112(.A1(358), .A2(18), .ZN(n176));
  XNOR2_X1  g0113(.A(n176), .B(n175), .ZN(n177));
  NOR2_X1   g0114(.A1(n133), .A2(n131), .ZN(n178));
  AOI21_X1  g0115(.A(n178), .B1(n136), .B2(n134), .ZN(n179));
  XOR2_X1   g0116(.A(n179), .B(n177), .ZN(n180));
  AND2_X1   g0117(.A1(375), .A2(\1 ), .ZN(n181));
  INV_X1    g0118(.A(n181), .ZN(n182));
  XNOR2_X1  g0119(.A(n182), .B(n180), .ZN(3211));
  AND4_X1   g0120(.A1(273), .A2(120), .A3(103), .A4(290), .ZN(n184));
  AOI22_X1  g0121(.A1(273), .A2(120), .B1(103), .B2(290), .ZN(n185));
  NOR2_X1   g0122(.A1(n185), .A2(n184), .ZN(n186));
  XNOR2_X1  g0123(.A(n186), .B(n138), .ZN(n187));
  AND2_X1   g0124(.A1(307), .A2(86), .ZN(n188));
  XNOR2_X1  g0125(.A(n188), .B(n187), .ZN(n189));
  NOR2_X1   g0126(.A1(n140), .A2(n105), .ZN(n190));
  OAI21_X1  g0127(.A(n105), .B1(n139), .B2(n138), .ZN(n191));
  OR3_X1    g0128(.A1(n139), .A2(n138), .A3(n105), .ZN(n192));
  AOI21_X1  g0129(.A(n142), .B1(n192), .B2(n191), .ZN(n193));
  NOR2_X1   g0130(.A1(n193), .A2(n190), .ZN(n194));
  XNOR2_X1  g0131(.A(n194), .B(n189), .ZN(n195));
  AND2_X1   g0132(.A1(324), .A2(69), .ZN(n196));
  XNOR2_X1  g0133(.A(n196), .B(n195), .ZN(n197));
  NOR2_X1   g0134(.A1(n148), .A2(n143), .ZN(n198));
  OR2_X1    g0135(.A1(n107), .A2(n85), .ZN(n199));
  NAND2_X1  g0136(.A1(307), .A2(69), .ZN(n200));
  AOI21_X1  g0137(.A(n200), .B1(n192), .B2(n191), .ZN(n201));
  AND3_X1   g0138(.A1(n200), .A2(n192), .A3(n191), .ZN(n202));
  OAI221_X1 g0139(.A(n199), .B1(n109), .B2(n108), .C1(n202), .C2(n201), .ZN(n203));
  NAND3_X1  g0140(.A1(n200), .A2(n192), .A3(n191), .ZN(n204));
  OAI221_X1 g0141(.A(n204), .B1(n141), .B2(n193), .C1(n147), .C2(n144), .ZN(n205));
  AOI21_X1  g0142(.A(n150), .B1(n205), .B2(n203), .ZN(n206));
  NOR2_X1   g0143(.A1(n206), .A2(n198), .ZN(n207));
  XNOR2_X1  g0144(.A(n207), .B(n197), .ZN(n208));
  AND2_X1   g0145(.A1(341), .A2(52), .ZN(n209));
  XNOR2_X1  g0146(.A(n209), .B(n208), .ZN(n210));
  NOR2_X1   g0147(.A1(n161), .A2(n151), .ZN(n211));
  OAI22_X1  g0148(.A1(n155), .A2(n156), .B1(n114), .B2(n111), .ZN(n212));
  INV_X1    g0149(.A(n150), .ZN(n213));
  AOI21_X1  g0150(.A(n213), .B1(n205), .B2(n203), .ZN(n214));
  AND3_X1   g0151(.A1(n213), .A2(n205), .A3(n203), .ZN(n215));
  OAI221_X1 g0152(.A(n212), .B1(n117), .B2(n116), .C1(n215), .C2(n214), .ZN(n216));
  NAND3_X1  g0153(.A1(n213), .A2(n205), .A3(n203), .ZN(n217));
  OAI221_X1 g0154(.A(n217), .B1(n149), .B2(n206), .C1(n160), .C2(n152), .ZN(n218));
  AOI21_X1  g0155(.A(n163), .B1(n218), .B2(n216), .ZN(n219));
  NOR2_X1   g0156(.A1(n219), .A2(n211), .ZN(n220));
  XNOR2_X1  g0157(.A(n220), .B(n210), .ZN(n221));
  AND2_X1   g0158(.A1(358), .A2(35), .ZN(n222));
  XNOR2_X1  g0159(.A(n222), .B(n221), .ZN(n223));
  NOR2_X1   g0160(.A1(n174), .A2(n164), .ZN(n224));
  OAI22_X1  g0161(.A1(n168), .A2(n169), .B1(n127), .B2(n119), .ZN(n225));
  INV_X1    g0162(.A(n163), .ZN(n226));
  AOI21_X1  g0163(.A(n226), .B1(n218), .B2(n216), .ZN(n227));
  AND3_X1   g0164(.A1(n226), .A2(n218), .A3(n216), .ZN(n228));
  OAI221_X1 g0165(.A(n225), .B1(n130), .B2(n129), .C1(n228), .C2(n227), .ZN(n229));
  NAND3_X1  g0166(.A1(n226), .A2(n218), .A3(n216), .ZN(n230));
  OAI221_X1 g0167(.A(n230), .B1(n162), .B2(n219), .C1(n173), .C2(n165), .ZN(n231));
  AOI21_X1  g0168(.A(n176), .B1(n231), .B2(n229), .ZN(n232));
  NOR2_X1   g0169(.A1(n232), .A2(n224), .ZN(n233));
  XNOR2_X1  g0170(.A(n233), .B(n223), .ZN(n234));
  AND2_X1   g0171(.A1(375), .A2(18), .ZN(n235));
  XNOR2_X1  g0172(.A(n235), .B(n234), .ZN(n236));
  NOR2_X1   g0173(.A1(n179), .A2(n177), .ZN(n237));
  AOI21_X1  g0174(.A(n237), .B1(n182), .B2(n180), .ZN(n238));
  XOR2_X1   g0175(.A(n238), .B(n236), .ZN(n239));
  AND2_X1   g0176(.A1(392), .A2(\1 ), .ZN(n240));
  INV_X1    g0177(.A(n240), .ZN(n241));
  XNOR2_X1  g0178(.A(n241), .B(n239), .ZN(3552));
  AND4_X1   g0179(.A1(273), .A2(137), .A3(120), .A4(290), .ZN(n243));
  AOI22_X1  g0180(.A1(273), .A2(137), .B1(120), .B2(290), .ZN(n244));
  NOR2_X1   g0181(.A1(n244), .A2(n243), .ZN(n245));
  XNOR2_X1  g0182(.A(n245), .B(n184), .ZN(n246));
  AND2_X1   g0183(.A1(307), .A2(103), .ZN(n247));
  XNOR2_X1  g0184(.A(n247), .B(n246), .ZN(n248));
  NOR2_X1   g0185(.A1(n186), .A2(n138), .ZN(n249));
  OAI21_X1  g0186(.A(n138), .B1(n185), .B2(n184), .ZN(n250));
  OR3_X1    g0187(.A1(n185), .A2(n184), .A3(n138), .ZN(n251));
  AOI21_X1  g0188(.A(n188), .B1(n251), .B2(n250), .ZN(n252));
  NOR2_X1   g0189(.A1(n252), .A2(n249), .ZN(n253));
  XNOR2_X1  g0190(.A(n253), .B(n248), .ZN(n254));
  AND2_X1   g0191(.A1(324), .A2(86), .ZN(n255));
  XNOR2_X1  g0192(.A(n255), .B(n254), .ZN(n256));
  NOR2_X1   g0193(.A1(n194), .A2(n189), .ZN(n257));
  OR2_X1    g0194(.A1(n140), .A2(n105), .ZN(n258));
  NAND2_X1  g0195(.A1(307), .A2(86), .ZN(n259));
  AOI21_X1  g0196(.A(n259), .B1(n251), .B2(n250), .ZN(n260));
  AND3_X1   g0197(.A1(n259), .A2(n251), .A3(n250), .ZN(n261));
  OAI221_X1 g0198(.A(n258), .B1(n142), .B2(n141), .C1(n261), .C2(n260), .ZN(n262));
  NAND3_X1  g0199(.A1(n259), .A2(n251), .A3(n250), .ZN(n263));
  OAI221_X1 g0200(.A(n263), .B1(n187), .B2(n252), .C1(n193), .C2(n190), .ZN(n264));
  AOI21_X1  g0201(.A(n196), .B1(n264), .B2(n262), .ZN(n265));
  NOR2_X1   g0202(.A1(n265), .A2(n257), .ZN(n266));
  XNOR2_X1  g0203(.A(n266), .B(n256), .ZN(n267));
  AND2_X1   g0204(.A1(341), .A2(69), .ZN(n268));
  XNOR2_X1  g0205(.A(n268), .B(n267), .ZN(n269));
  NOR2_X1   g0206(.A1(n207), .A2(n197), .ZN(n270));
  OAI22_X1  g0207(.A1(n201), .A2(n202), .B1(n147), .B2(n144), .ZN(n271));
  INV_X1    g0208(.A(n196), .ZN(n272));
  AOI21_X1  g0209(.A(n272), .B1(n264), .B2(n262), .ZN(n273));
  AND3_X1   g0210(.A1(n272), .A2(n264), .A3(n262), .ZN(n274));
  OAI221_X1 g0211(.A(n271), .B1(n150), .B2(n149), .C1(n274), .C2(n273), .ZN(n275));
  NAND3_X1  g0212(.A1(n272), .A2(n264), .A3(n262), .ZN(n276));
  OAI221_X1 g0213(.A(n276), .B1(n195), .B2(n265), .C1(n206), .C2(n198), .ZN(n277));
  AOI21_X1  g0214(.A(n209), .B1(n277), .B2(n275), .ZN(n278));
  NOR2_X1   g0215(.A1(n278), .A2(n270), .ZN(n279));
  XNOR2_X1  g0216(.A(n279), .B(n269), .ZN(n280));
  AND2_X1   g0217(.A1(358), .A2(52), .ZN(n281));
  XNOR2_X1  g0218(.A(n281), .B(n280), .ZN(n282));
  NOR2_X1   g0219(.A1(n220), .A2(n210), .ZN(n283));
  OAI22_X1  g0220(.A1(n214), .A2(n215), .B1(n160), .B2(n152), .ZN(n284));
  INV_X1    g0221(.A(n209), .ZN(n285));
  AOI21_X1  g0222(.A(n285), .B1(n277), .B2(n275), .ZN(n286));
  AND3_X1   g0223(.A1(n285), .A2(n277), .A3(n275), .ZN(n287));
  OAI221_X1 g0224(.A(n284), .B1(n163), .B2(n162), .C1(n287), .C2(n286), .ZN(n288));
  NAND3_X1  g0225(.A1(n285), .A2(n277), .A3(n275), .ZN(n289));
  OAI221_X1 g0226(.A(n289), .B1(n208), .B2(n278), .C1(n219), .C2(n211), .ZN(n290));
  AOI21_X1  g0227(.A(n222), .B1(n290), .B2(n288), .ZN(n291));
  NOR2_X1   g0228(.A1(n291), .A2(n283), .ZN(n292));
  XNOR2_X1  g0229(.A(n292), .B(n282), .ZN(n293));
  AND2_X1   g0230(.A1(375), .A2(35), .ZN(n294));
  XNOR2_X1  g0231(.A(n294), .B(n293), .ZN(n295));
  NOR2_X1   g0232(.A1(n233), .A2(n223), .ZN(n296));
  OAI22_X1  g0233(.A1(n227), .A2(n228), .B1(n173), .B2(n165), .ZN(n297));
  INV_X1    g0234(.A(n222), .ZN(n298));
  AOI21_X1  g0235(.A(n298), .B1(n290), .B2(n288), .ZN(n299));
  AND3_X1   g0236(.A1(n298), .A2(n290), .A3(n288), .ZN(n300));
  OAI221_X1 g0237(.A(n297), .B1(n176), .B2(n175), .C1(n300), .C2(n299), .ZN(n301));
  NAND3_X1  g0238(.A1(n298), .A2(n290), .A3(n288), .ZN(n302));
  OAI221_X1 g0239(.A(n302), .B1(n221), .B2(n291), .C1(n232), .C2(n224), .ZN(n303));
  AOI21_X1  g0240(.A(n235), .B1(n303), .B2(n301), .ZN(n304));
  NOR2_X1   g0241(.A1(n304), .A2(n296), .ZN(n305));
  XNOR2_X1  g0242(.A(n305), .B(n295), .ZN(n306));
  AND2_X1   g0243(.A1(392), .A2(18), .ZN(n307));
  XNOR2_X1  g0244(.A(n307), .B(n306), .ZN(n308));
  NOR2_X1   g0245(.A1(n238), .A2(n236), .ZN(n309));
  AOI21_X1  g0246(.A(n309), .B1(n241), .B2(n239), .ZN(n310));
  XOR2_X1   g0247(.A(n310), .B(n308), .ZN(n311));
  AND2_X1   g0248(.A1(409), .A2(\1 ), .ZN(n312));
  INV_X1    g0249(.A(n312), .ZN(n313));
  XNOR2_X1  g0250(.A(n313), .B(n311), .ZN(3895));
  AND4_X1   g0251(.A1(273), .A2(154), .A3(137), .A4(290), .ZN(n315));
  AOI22_X1  g0252(.A1(273), .A2(154), .B1(137), .B2(290), .ZN(n316));
  NOR2_X1   g0253(.A1(n316), .A2(n315), .ZN(n317));
  XNOR2_X1  g0254(.A(n317), .B(n243), .ZN(n318));
  AND2_X1   g0255(.A1(307), .A2(120), .ZN(n319));
  XNOR2_X1  g0256(.A(n319), .B(n318), .ZN(n320));
  NOR2_X1   g0257(.A1(n245), .A2(n184), .ZN(n321));
  OAI21_X1  g0258(.A(n184), .B1(n244), .B2(n243), .ZN(n322));
  OR3_X1    g0259(.A1(n244), .A2(n243), .A3(n184), .ZN(n323));
  AOI21_X1  g0260(.A(n247), .B1(n323), .B2(n322), .ZN(n324));
  NOR2_X1   g0261(.A1(n324), .A2(n321), .ZN(n325));
  XNOR2_X1  g0262(.A(n325), .B(n320), .ZN(n326));
  AND2_X1   g0263(.A1(324), .A2(103), .ZN(n327));
  XNOR2_X1  g0264(.A(n327), .B(n326), .ZN(n328));
  NOR2_X1   g0265(.A1(n253), .A2(n248), .ZN(n329));
  OR2_X1    g0266(.A1(n186), .A2(n138), .ZN(n330));
  NAND2_X1  g0267(.A1(307), .A2(103), .ZN(n331));
  AOI21_X1  g0268(.A(n331), .B1(n323), .B2(n322), .ZN(n332));
  AND3_X1   g0269(.A1(n331), .A2(n323), .A3(n322), .ZN(n333));
  OAI221_X1 g0270(.A(n330), .B1(n188), .B2(n187), .C1(n333), .C2(n332), .ZN(n334));
  NAND3_X1  g0271(.A1(n331), .A2(n323), .A3(n322), .ZN(n335));
  OAI221_X1 g0272(.A(n335), .B1(n246), .B2(n324), .C1(n252), .C2(n249), .ZN(n336));
  AOI21_X1  g0273(.A(n255), .B1(n336), .B2(n334), .ZN(n337));
  NOR2_X1   g0274(.A1(n337), .A2(n329), .ZN(n338));
  XNOR2_X1  g0275(.A(n338), .B(n328), .ZN(n339));
  AND2_X1   g0276(.A1(341), .A2(86), .ZN(n340));
  XNOR2_X1  g0277(.A(n340), .B(n339), .ZN(n341));
  NOR2_X1   g0278(.A1(n266), .A2(n256), .ZN(n342));
  OAI22_X1  g0279(.A1(n260), .A2(n261), .B1(n193), .B2(n190), .ZN(n343));
  INV_X1    g0280(.A(n255), .ZN(n344));
  AOI21_X1  g0281(.A(n344), .B1(n336), .B2(n334), .ZN(n345));
  AND3_X1   g0282(.A1(n344), .A2(n336), .A3(n334), .ZN(n346));
  OAI221_X1 g0283(.A(n343), .B1(n196), .B2(n195), .C1(n346), .C2(n345), .ZN(n347));
  NAND3_X1  g0284(.A1(n344), .A2(n336), .A3(n334), .ZN(n348));
  OAI221_X1 g0285(.A(n348), .B1(n254), .B2(n337), .C1(n265), .C2(n257), .ZN(n349));
  AOI21_X1  g0286(.A(n268), .B1(n349), .B2(n347), .ZN(n350));
  NOR2_X1   g0287(.A1(n350), .A2(n342), .ZN(n351));
  XNOR2_X1  g0288(.A(n351), .B(n341), .ZN(n352));
  AND2_X1   g0289(.A1(358), .A2(69), .ZN(n353));
  XNOR2_X1  g0290(.A(n353), .B(n352), .ZN(n354));
  NOR2_X1   g0291(.A1(n279), .A2(n269), .ZN(n355));
  OAI22_X1  g0292(.A1(n273), .A2(n274), .B1(n206), .B2(n198), .ZN(n356));
  INV_X1    g0293(.A(n268), .ZN(n357));
  AOI21_X1  g0294(.A(n357), .B1(n349), .B2(n347), .ZN(n358));
  AND3_X1   g0295(.A1(n357), .A2(n349), .A3(n347), .ZN(n359));
  OAI221_X1 g0296(.A(n356), .B1(n209), .B2(n208), .C1(n359), .C2(n358), .ZN(n360));
  NAND3_X1  g0297(.A1(n357), .A2(n349), .A3(n347), .ZN(n361));
  OAI221_X1 g0298(.A(n361), .B1(n267), .B2(n350), .C1(n278), .C2(n270), .ZN(n362));
  AOI21_X1  g0299(.A(n281), .B1(n362), .B2(n360), .ZN(n363));
  NOR2_X1   g0300(.A1(n363), .A2(n355), .ZN(n364));
  XNOR2_X1  g0301(.A(n364), .B(n354), .ZN(n365));
  AND2_X1   g0302(.A1(375), .A2(52), .ZN(n366));
  XNOR2_X1  g0303(.A(n366), .B(n365), .ZN(n367));
  NOR2_X1   g0304(.A1(n292), .A2(n282), .ZN(n368));
  OAI22_X1  g0305(.A1(n286), .A2(n287), .B1(n219), .B2(n211), .ZN(n369));
  INV_X1    g0306(.A(n281), .ZN(n370));
  AOI21_X1  g0307(.A(n370), .B1(n362), .B2(n360), .ZN(n371));
  AND3_X1   g0308(.A1(n370), .A2(n362), .A3(n360), .ZN(n372));
  OAI221_X1 g0309(.A(n369), .B1(n222), .B2(n221), .C1(n372), .C2(n371), .ZN(n373));
  NAND3_X1  g0310(.A1(n370), .A2(n362), .A3(n360), .ZN(n374));
  OAI221_X1 g0311(.A(n374), .B1(n280), .B2(n363), .C1(n291), .C2(n283), .ZN(n375));
  AOI21_X1  g0312(.A(n294), .B1(n375), .B2(n373), .ZN(n376));
  NOR2_X1   g0313(.A1(n376), .A2(n368), .ZN(n377));
  XNOR2_X1  g0314(.A(n377), .B(n367), .ZN(n378));
  AND2_X1   g0315(.A1(392), .A2(35), .ZN(n379));
  XNOR2_X1  g0316(.A(n379), .B(n378), .ZN(n380));
  NOR2_X1   g0317(.A1(n305), .A2(n295), .ZN(n381));
  OAI22_X1  g0318(.A1(n299), .A2(n300), .B1(n232), .B2(n224), .ZN(n382));
  INV_X1    g0319(.A(n294), .ZN(n383));
  AOI21_X1  g0320(.A(n383), .B1(n375), .B2(n373), .ZN(n384));
  AND3_X1   g0321(.A1(n383), .A2(n375), .A3(n373), .ZN(n385));
  OAI221_X1 g0322(.A(n382), .B1(n235), .B2(n234), .C1(n385), .C2(n384), .ZN(n386));
  NAND3_X1  g0323(.A1(n383), .A2(n375), .A3(n373), .ZN(n387));
  OAI221_X1 g0324(.A(n387), .B1(n293), .B2(n376), .C1(n304), .C2(n296), .ZN(n388));
  AOI21_X1  g0325(.A(n307), .B1(n388), .B2(n386), .ZN(n389));
  NOR2_X1   g0326(.A1(n389), .A2(n381), .ZN(n390));
  XNOR2_X1  g0327(.A(n390), .B(n380), .ZN(n391));
  AND2_X1   g0328(.A1(409), .A2(18), .ZN(n392));
  XNOR2_X1  g0329(.A(n392), .B(n391), .ZN(n393));
  NOR2_X1   g0330(.A1(n310), .A2(n308), .ZN(n394));
  AOI21_X1  g0331(.A(n394), .B1(n313), .B2(n311), .ZN(n395));
  XOR2_X1   g0332(.A(n395), .B(n393), .ZN(n396));
  AND2_X1   g0333(.A1(426), .A2(\1 ), .ZN(n397));
  INV_X1    g0334(.A(n397), .ZN(n398));
  XNOR2_X1  g0335(.A(n398), .B(n396), .ZN(4241));
  AND4_X1   g0336(.A1(273), .A2(171), .A3(154), .A4(290), .ZN(n400));
  AOI22_X1  g0337(.A1(273), .A2(171), .B1(154), .B2(290), .ZN(n401));
  NOR2_X1   g0338(.A1(n401), .A2(n400), .ZN(n402));
  XNOR2_X1  g0339(.A(n402), .B(n315), .ZN(n403));
  AND2_X1   g0340(.A1(307), .A2(137), .ZN(n404));
  XNOR2_X1  g0341(.A(n404), .B(n403), .ZN(n405));
  NOR2_X1   g0342(.A1(n317), .A2(n243), .ZN(n406));
  OAI21_X1  g0343(.A(n243), .B1(n316), .B2(n315), .ZN(n407));
  OR3_X1    g0344(.A1(n316), .A2(n315), .A3(n243), .ZN(n408));
  AOI21_X1  g0345(.A(n319), .B1(n408), .B2(n407), .ZN(n409));
  NOR2_X1   g0346(.A1(n409), .A2(n406), .ZN(n410));
  XNOR2_X1  g0347(.A(n410), .B(n405), .ZN(n411));
  AND2_X1   g0348(.A1(324), .A2(120), .ZN(n412));
  XNOR2_X1  g0349(.A(n412), .B(n411), .ZN(n413));
  NOR2_X1   g0350(.A1(n325), .A2(n320), .ZN(n414));
  OR2_X1    g0351(.A1(n245), .A2(n184), .ZN(n415));
  NAND2_X1  g0352(.A1(307), .A2(120), .ZN(n416));
  AOI21_X1  g0353(.A(n416), .B1(n408), .B2(n407), .ZN(n417));
  AND3_X1   g0354(.A1(n416), .A2(n408), .A3(n407), .ZN(n418));
  OAI221_X1 g0355(.A(n415), .B1(n247), .B2(n246), .C1(n418), .C2(n417), .ZN(n419));
  NAND3_X1  g0356(.A1(n416), .A2(n408), .A3(n407), .ZN(n420));
  OAI221_X1 g0357(.A(n420), .B1(n318), .B2(n409), .C1(n324), .C2(n321), .ZN(n421));
  AOI21_X1  g0358(.A(n327), .B1(n421), .B2(n419), .ZN(n422));
  NOR2_X1   g0359(.A1(n422), .A2(n414), .ZN(n423));
  XNOR2_X1  g0360(.A(n423), .B(n413), .ZN(n424));
  AND2_X1   g0361(.A1(341), .A2(103), .ZN(n425));
  XNOR2_X1  g0362(.A(n425), .B(n424), .ZN(n426));
  NOR2_X1   g0363(.A1(n338), .A2(n328), .ZN(n427));
  OAI22_X1  g0364(.A1(n332), .A2(n333), .B1(n252), .B2(n249), .ZN(n428));
  INV_X1    g0365(.A(n327), .ZN(n429));
  AOI21_X1  g0366(.A(n429), .B1(n421), .B2(n419), .ZN(n430));
  AND3_X1   g0367(.A1(n429), .A2(n421), .A3(n419), .ZN(n431));
  OAI221_X1 g0368(.A(n428), .B1(n255), .B2(n254), .C1(n431), .C2(n430), .ZN(n432));
  NAND3_X1  g0369(.A1(n429), .A2(n421), .A3(n419), .ZN(n433));
  OAI221_X1 g0370(.A(n433), .B1(n326), .B2(n422), .C1(n337), .C2(n329), .ZN(n434));
  AOI21_X1  g0371(.A(n340), .B1(n434), .B2(n432), .ZN(n435));
  NOR2_X1   g0372(.A1(n435), .A2(n427), .ZN(n436));
  XNOR2_X1  g0373(.A(n436), .B(n426), .ZN(n437));
  AND2_X1   g0374(.A1(358), .A2(86), .ZN(n438));
  XNOR2_X1  g0375(.A(n438), .B(n437), .ZN(n439));
  NOR2_X1   g0376(.A1(n351), .A2(n341), .ZN(n440));
  OAI22_X1  g0377(.A1(n345), .A2(n346), .B1(n265), .B2(n257), .ZN(n441));
  INV_X1    g0378(.A(n340), .ZN(n442));
  AOI21_X1  g0379(.A(n442), .B1(n434), .B2(n432), .ZN(n443));
  AND3_X1   g0380(.A1(n442), .A2(n434), .A3(n432), .ZN(n444));
  OAI221_X1 g0381(.A(n441), .B1(n268), .B2(n267), .C1(n444), .C2(n443), .ZN(n445));
  NAND3_X1  g0382(.A1(n442), .A2(n434), .A3(n432), .ZN(n446));
  OAI221_X1 g0383(.A(n446), .B1(n339), .B2(n435), .C1(n350), .C2(n342), .ZN(n447));
  AOI21_X1  g0384(.A(n353), .B1(n447), .B2(n445), .ZN(n448));
  NOR2_X1   g0385(.A1(n448), .A2(n440), .ZN(n449));
  XNOR2_X1  g0386(.A(n449), .B(n439), .ZN(n450));
  AND2_X1   g0387(.A1(375), .A2(69), .ZN(n451));
  XNOR2_X1  g0388(.A(n451), .B(n450), .ZN(n452));
  NOR2_X1   g0389(.A1(n364), .A2(n354), .ZN(n453));
  OAI22_X1  g0390(.A1(n358), .A2(n359), .B1(n278), .B2(n270), .ZN(n454));
  INV_X1    g0391(.A(n353), .ZN(n455));
  AOI21_X1  g0392(.A(n455), .B1(n447), .B2(n445), .ZN(n456));
  AND3_X1   g0393(.A1(n455), .A2(n447), .A3(n445), .ZN(n457));
  OAI221_X1 g0394(.A(n454), .B1(n281), .B2(n280), .C1(n457), .C2(n456), .ZN(n458));
  NAND3_X1  g0395(.A1(n455), .A2(n447), .A3(n445), .ZN(n459));
  OAI221_X1 g0396(.A(n459), .B1(n352), .B2(n448), .C1(n363), .C2(n355), .ZN(n460));
  AOI21_X1  g0397(.A(n366), .B1(n460), .B2(n458), .ZN(n461));
  NOR2_X1   g0398(.A1(n461), .A2(n453), .ZN(n462));
  XNOR2_X1  g0399(.A(n462), .B(n452), .ZN(n463));
  AND2_X1   g0400(.A1(392), .A2(52), .ZN(n464));
  XNOR2_X1  g0401(.A(n464), .B(n463), .ZN(n465));
  NOR2_X1   g0402(.A1(n377), .A2(n367), .ZN(n466));
  OAI22_X1  g0403(.A1(n371), .A2(n372), .B1(n291), .B2(n283), .ZN(n467));
  INV_X1    g0404(.A(n366), .ZN(n468));
  AOI21_X1  g0405(.A(n468), .B1(n460), .B2(n458), .ZN(n469));
  AND3_X1   g0406(.A1(n468), .A2(n460), .A3(n458), .ZN(n470));
  OAI221_X1 g0407(.A(n467), .B1(n294), .B2(n293), .C1(n470), .C2(n469), .ZN(n471));
  NAND3_X1  g0408(.A1(n468), .A2(n460), .A3(n458), .ZN(n472));
  OAI221_X1 g0409(.A(n472), .B1(n365), .B2(n461), .C1(n376), .C2(n368), .ZN(n473));
  AOI21_X1  g0410(.A(n379), .B1(n473), .B2(n471), .ZN(n474));
  NOR2_X1   g0411(.A1(n474), .A2(n466), .ZN(n475));
  XNOR2_X1  g0412(.A(n475), .B(n465), .ZN(n476));
  AND2_X1   g0413(.A1(409), .A2(35), .ZN(n477));
  XNOR2_X1  g0414(.A(n477), .B(n476), .ZN(n478));
  NOR2_X1   g0415(.A1(n390), .A2(n380), .ZN(n479));
  OAI22_X1  g0416(.A1(n384), .A2(n385), .B1(n304), .B2(n296), .ZN(n480));
  INV_X1    g0417(.A(n379), .ZN(n481));
  AOI21_X1  g0418(.A(n481), .B1(n473), .B2(n471), .ZN(n482));
  AND3_X1   g0419(.A1(n481), .A2(n473), .A3(n471), .ZN(n483));
  OAI221_X1 g0420(.A(n480), .B1(n307), .B2(n306), .C1(n483), .C2(n482), .ZN(n484));
  NAND3_X1  g0421(.A1(n481), .A2(n473), .A3(n471), .ZN(n485));
  OAI221_X1 g0422(.A(n485), .B1(n378), .B2(n474), .C1(n389), .C2(n381), .ZN(n486));
  AOI21_X1  g0423(.A(n392), .B1(n486), .B2(n484), .ZN(n487));
  NOR2_X1   g0424(.A1(n487), .A2(n479), .ZN(n488));
  XNOR2_X1  g0425(.A(n488), .B(n478), .ZN(n489));
  AND2_X1   g0426(.A1(426), .A2(18), .ZN(n490));
  XNOR2_X1  g0427(.A(n490), .B(n489), .ZN(n491));
  NOR2_X1   g0428(.A1(n395), .A2(n393), .ZN(n492));
  AOI21_X1  g0429(.A(n492), .B1(n398), .B2(n396), .ZN(n493));
  XOR2_X1   g0430(.A(n493), .B(n491), .ZN(n494));
  AND2_X1   g0431(.A1(443), .A2(\1 ), .ZN(n495));
  INV_X1    g0432(.A(n495), .ZN(n496));
  XNOR2_X1  g0433(.A(n496), .B(n494), .ZN(4591));
  AND4_X1   g0434(.A1(273), .A2(188), .A3(171), .A4(290), .ZN(n498));
  AOI22_X1  g0435(.A1(273), .A2(188), .B1(171), .B2(290), .ZN(n499));
  NOR2_X1   g0436(.A1(n499), .A2(n498), .ZN(n500));
  XNOR2_X1  g0437(.A(n500), .B(n400), .ZN(n501));
  AND2_X1   g0438(.A1(307), .A2(154), .ZN(n502));
  XNOR2_X1  g0439(.A(n502), .B(n501), .ZN(n503));
  NOR2_X1   g0440(.A1(n402), .A2(n315), .ZN(n504));
  OAI21_X1  g0441(.A(n315), .B1(n401), .B2(n400), .ZN(n505));
  OR3_X1    g0442(.A1(n401), .A2(n400), .A3(n315), .ZN(n506));
  AOI21_X1  g0443(.A(n404), .B1(n506), .B2(n505), .ZN(n507));
  NOR2_X1   g0444(.A1(n507), .A2(n504), .ZN(n508));
  XNOR2_X1  g0445(.A(n508), .B(n503), .ZN(n509));
  AND2_X1   g0446(.A1(324), .A2(137), .ZN(n510));
  XNOR2_X1  g0447(.A(n510), .B(n509), .ZN(n511));
  NOR2_X1   g0448(.A1(n410), .A2(n405), .ZN(n512));
  OR2_X1    g0449(.A1(n317), .A2(n243), .ZN(n513));
  NAND2_X1  g0450(.A1(307), .A2(137), .ZN(n514));
  AOI21_X1  g0451(.A(n514), .B1(n506), .B2(n505), .ZN(n515));
  AND3_X1   g0452(.A1(n514), .A2(n506), .A3(n505), .ZN(n516));
  OAI221_X1 g0453(.A(n513), .B1(n319), .B2(n318), .C1(n516), .C2(n515), .ZN(n517));
  NAND3_X1  g0454(.A1(n514), .A2(n506), .A3(n505), .ZN(n518));
  OAI221_X1 g0455(.A(n518), .B1(n403), .B2(n507), .C1(n409), .C2(n406), .ZN(n519));
  AOI21_X1  g0456(.A(n412), .B1(n519), .B2(n517), .ZN(n520));
  NOR2_X1   g0457(.A1(n520), .A2(n512), .ZN(n521));
  XNOR2_X1  g0458(.A(n521), .B(n511), .ZN(n522));
  AND2_X1   g0459(.A1(341), .A2(120), .ZN(n523));
  XNOR2_X1  g0460(.A(n523), .B(n522), .ZN(n524));
  NOR2_X1   g0461(.A1(n423), .A2(n413), .ZN(n525));
  OAI22_X1  g0462(.A1(n417), .A2(n418), .B1(n324), .B2(n321), .ZN(n526));
  INV_X1    g0463(.A(n412), .ZN(n527));
  AOI21_X1  g0464(.A(n527), .B1(n519), .B2(n517), .ZN(n528));
  AND3_X1   g0465(.A1(n527), .A2(n519), .A3(n517), .ZN(n529));
  OAI221_X1 g0466(.A(n526), .B1(n327), .B2(n326), .C1(n529), .C2(n528), .ZN(n530));
  NAND3_X1  g0467(.A1(n527), .A2(n519), .A3(n517), .ZN(n531));
  OAI221_X1 g0468(.A(n531), .B1(n411), .B2(n520), .C1(n422), .C2(n414), .ZN(n532));
  AOI21_X1  g0469(.A(n425), .B1(n532), .B2(n530), .ZN(n533));
  NOR2_X1   g0470(.A1(n533), .A2(n525), .ZN(n534));
  XNOR2_X1  g0471(.A(n534), .B(n524), .ZN(n535));
  AND2_X1   g0472(.A1(358), .A2(103), .ZN(n536));
  XNOR2_X1  g0473(.A(n536), .B(n535), .ZN(n537));
  NOR2_X1   g0474(.A1(n436), .A2(n426), .ZN(n538));
  OAI22_X1  g0475(.A1(n430), .A2(n431), .B1(n337), .B2(n329), .ZN(n539));
  INV_X1    g0476(.A(n425), .ZN(n540));
  AOI21_X1  g0477(.A(n540), .B1(n532), .B2(n530), .ZN(n541));
  AND3_X1   g0478(.A1(n540), .A2(n532), .A3(n530), .ZN(n542));
  OAI221_X1 g0479(.A(n539), .B1(n340), .B2(n339), .C1(n542), .C2(n541), .ZN(n543));
  NAND3_X1  g0480(.A1(n540), .A2(n532), .A3(n530), .ZN(n544));
  OAI221_X1 g0481(.A(n544), .B1(n424), .B2(n533), .C1(n435), .C2(n427), .ZN(n545));
  AOI21_X1  g0482(.A(n438), .B1(n545), .B2(n543), .ZN(n546));
  NOR2_X1   g0483(.A1(n546), .A2(n538), .ZN(n547));
  XNOR2_X1  g0484(.A(n547), .B(n537), .ZN(n548));
  AND2_X1   g0485(.A1(375), .A2(86), .ZN(n549));
  XNOR2_X1  g0486(.A(n549), .B(n548), .ZN(n550));
  NOR2_X1   g0487(.A1(n449), .A2(n439), .ZN(n551));
  OAI22_X1  g0488(.A1(n443), .A2(n444), .B1(n350), .B2(n342), .ZN(n552));
  INV_X1    g0489(.A(n438), .ZN(n553));
  AOI21_X1  g0490(.A(n553), .B1(n545), .B2(n543), .ZN(n554));
  AND3_X1   g0491(.A1(n553), .A2(n545), .A3(n543), .ZN(n555));
  OAI221_X1 g0492(.A(n552), .B1(n353), .B2(n352), .C1(n555), .C2(n554), .ZN(n556));
  NAND3_X1  g0493(.A1(n553), .A2(n545), .A3(n543), .ZN(n557));
  OAI221_X1 g0494(.A(n557), .B1(n437), .B2(n546), .C1(n448), .C2(n440), .ZN(n558));
  AOI21_X1  g0495(.A(n451), .B1(n558), .B2(n556), .ZN(n559));
  NOR2_X1   g0496(.A1(n559), .A2(n551), .ZN(n560));
  XNOR2_X1  g0497(.A(n560), .B(n550), .ZN(n561));
  AND2_X1   g0498(.A1(392), .A2(69), .ZN(n562));
  XNOR2_X1  g0499(.A(n562), .B(n561), .ZN(n563));
  NOR2_X1   g0500(.A1(n462), .A2(n452), .ZN(n564));
  OAI22_X1  g0501(.A1(n456), .A2(n457), .B1(n363), .B2(n355), .ZN(n565));
  INV_X1    g0502(.A(n451), .ZN(n566));
  AOI21_X1  g0503(.A(n566), .B1(n558), .B2(n556), .ZN(n567));
  AND3_X1   g0504(.A1(n566), .A2(n558), .A3(n556), .ZN(n568));
  OAI221_X1 g0505(.A(n565), .B1(n366), .B2(n365), .C1(n568), .C2(n567), .ZN(n569));
  NAND3_X1  g0506(.A1(n566), .A2(n558), .A3(n556), .ZN(n570));
  OAI221_X1 g0507(.A(n570), .B1(n450), .B2(n559), .C1(n461), .C2(n453), .ZN(n571));
  AOI21_X1  g0508(.A(n464), .B1(n571), .B2(n569), .ZN(n572));
  NOR2_X1   g0509(.A1(n572), .A2(n564), .ZN(n573));
  XNOR2_X1  g0510(.A(n573), .B(n563), .ZN(n574));
  AND2_X1   g0511(.A1(409), .A2(52), .ZN(n575));
  XNOR2_X1  g0512(.A(n575), .B(n574), .ZN(n576));
  NOR2_X1   g0513(.A1(n475), .A2(n465), .ZN(n577));
  OAI22_X1  g0514(.A1(n469), .A2(n470), .B1(n376), .B2(n368), .ZN(n578));
  INV_X1    g0515(.A(n464), .ZN(n579));
  AOI21_X1  g0516(.A(n579), .B1(n571), .B2(n569), .ZN(n580));
  AND3_X1   g0517(.A1(n579), .A2(n571), .A3(n569), .ZN(n581));
  OAI221_X1 g0518(.A(n578), .B1(n379), .B2(n378), .C1(n581), .C2(n580), .ZN(n582));
  NAND3_X1  g0519(.A1(n579), .A2(n571), .A3(n569), .ZN(n583));
  OAI221_X1 g0520(.A(n583), .B1(n463), .B2(n572), .C1(n474), .C2(n466), .ZN(n584));
  AOI21_X1  g0521(.A(n477), .B1(n584), .B2(n582), .ZN(n585));
  NOR2_X1   g0522(.A1(n585), .A2(n577), .ZN(n586));
  XNOR2_X1  g0523(.A(n586), .B(n576), .ZN(n587));
  AND2_X1   g0524(.A1(426), .A2(35), .ZN(n588));
  XNOR2_X1  g0525(.A(n588), .B(n587), .ZN(n589));
  NOR2_X1   g0526(.A1(n488), .A2(n478), .ZN(n590));
  OAI22_X1  g0527(.A1(n482), .A2(n483), .B1(n389), .B2(n381), .ZN(n591));
  INV_X1    g0528(.A(n477), .ZN(n592));
  AOI21_X1  g0529(.A(n592), .B1(n584), .B2(n582), .ZN(n593));
  AND3_X1   g0530(.A1(n592), .A2(n584), .A3(n582), .ZN(n594));
  OAI221_X1 g0531(.A(n591), .B1(n392), .B2(n391), .C1(n594), .C2(n593), .ZN(n595));
  NAND3_X1  g0532(.A1(n592), .A2(n584), .A3(n582), .ZN(n596));
  OAI221_X1 g0533(.A(n596), .B1(n476), .B2(n585), .C1(n487), .C2(n479), .ZN(n597));
  AOI21_X1  g0534(.A(n490), .B1(n597), .B2(n595), .ZN(n598));
  NOR2_X1   g0535(.A1(n598), .A2(n590), .ZN(n599));
  XNOR2_X1  g0536(.A(n599), .B(n589), .ZN(n600));
  AND2_X1   g0537(.A1(443), .A2(18), .ZN(n601));
  XNOR2_X1  g0538(.A(n601), .B(n600), .ZN(n602));
  NOR2_X1   g0539(.A1(n493), .A2(n491), .ZN(n603));
  AOI21_X1  g0540(.A(n603), .B1(n496), .B2(n494), .ZN(n604));
  XOR2_X1   g0541(.A(n604), .B(n602), .ZN(n605));
  AND2_X1   g0542(.A1(460), .A2(\1 ), .ZN(n606));
  INV_X1    g0543(.A(n606), .ZN(n607));
  XNOR2_X1  g0544(.A(n607), .B(n605), .ZN(4946));
  AND4_X1   g0545(.A1(273), .A2(205), .A3(188), .A4(290), .ZN(n609));
  AOI22_X1  g0546(.A1(273), .A2(205), .B1(188), .B2(290), .ZN(n610));
  NOR2_X1   g0547(.A1(n610), .A2(n609), .ZN(n611));
  XNOR2_X1  g0548(.A(n611), .B(n498), .ZN(n612));
  AND2_X1   g0549(.A1(307), .A2(171), .ZN(n613));
  XNOR2_X1  g0550(.A(n613), .B(n612), .ZN(n614));
  NOR2_X1   g0551(.A1(n500), .A2(n400), .ZN(n615));
  OAI21_X1  g0552(.A(n400), .B1(n499), .B2(n498), .ZN(n616));
  OR3_X1    g0553(.A1(n499), .A2(n498), .A3(n400), .ZN(n617));
  AOI21_X1  g0554(.A(n502), .B1(n617), .B2(n616), .ZN(n618));
  NOR2_X1   g0555(.A1(n618), .A2(n615), .ZN(n619));
  XNOR2_X1  g0556(.A(n619), .B(n614), .ZN(n620));
  AND2_X1   g0557(.A1(324), .A2(154), .ZN(n621));
  XNOR2_X1  g0558(.A(n621), .B(n620), .ZN(n622));
  NOR2_X1   g0559(.A1(n508), .A2(n503), .ZN(n623));
  OR2_X1    g0560(.A1(n402), .A2(n315), .ZN(n624));
  NAND2_X1  g0561(.A1(307), .A2(154), .ZN(n625));
  AOI21_X1  g0562(.A(n625), .B1(n617), .B2(n616), .ZN(n626));
  AND3_X1   g0563(.A1(n625), .A2(n617), .A3(n616), .ZN(n627));
  OAI221_X1 g0564(.A(n624), .B1(n404), .B2(n403), .C1(n627), .C2(n626), .ZN(n628));
  NAND3_X1  g0565(.A1(n625), .A2(n617), .A3(n616), .ZN(n629));
  OAI221_X1 g0566(.A(n629), .B1(n501), .B2(n618), .C1(n507), .C2(n504), .ZN(n630));
  AOI21_X1  g0567(.A(n510), .B1(n630), .B2(n628), .ZN(n631));
  NOR2_X1   g0568(.A1(n631), .A2(n623), .ZN(n632));
  XNOR2_X1  g0569(.A(n632), .B(n622), .ZN(n633));
  AND2_X1   g0570(.A1(341), .A2(137), .ZN(n634));
  XNOR2_X1  g0571(.A(n634), .B(n633), .ZN(n635));
  NOR2_X1   g0572(.A1(n521), .A2(n511), .ZN(n636));
  OAI22_X1  g0573(.A1(n515), .A2(n516), .B1(n409), .B2(n406), .ZN(n637));
  INV_X1    g0574(.A(n510), .ZN(n638));
  AOI21_X1  g0575(.A(n638), .B1(n630), .B2(n628), .ZN(n639));
  AND3_X1   g0576(.A1(n638), .A2(n630), .A3(n628), .ZN(n640));
  OAI221_X1 g0577(.A(n637), .B1(n412), .B2(n411), .C1(n640), .C2(n639), .ZN(n641));
  NAND3_X1  g0578(.A1(n638), .A2(n630), .A3(n628), .ZN(n642));
  OAI221_X1 g0579(.A(n642), .B1(n509), .B2(n631), .C1(n520), .C2(n512), .ZN(n643));
  AOI21_X1  g0580(.A(n523), .B1(n643), .B2(n641), .ZN(n644));
  NOR2_X1   g0581(.A1(n644), .A2(n636), .ZN(n645));
  XNOR2_X1  g0582(.A(n645), .B(n635), .ZN(n646));
  AND2_X1   g0583(.A1(358), .A2(120), .ZN(n647));
  XNOR2_X1  g0584(.A(n647), .B(n646), .ZN(n648));
  NOR2_X1   g0585(.A1(n534), .A2(n524), .ZN(n649));
  OAI22_X1  g0586(.A1(n528), .A2(n529), .B1(n422), .B2(n414), .ZN(n650));
  INV_X1    g0587(.A(n523), .ZN(n651));
  AOI21_X1  g0588(.A(n651), .B1(n643), .B2(n641), .ZN(n652));
  AND3_X1   g0589(.A1(n651), .A2(n643), .A3(n641), .ZN(n653));
  OAI221_X1 g0590(.A(n650), .B1(n425), .B2(n424), .C1(n653), .C2(n652), .ZN(n654));
  NAND3_X1  g0591(.A1(n651), .A2(n643), .A3(n641), .ZN(n655));
  OAI221_X1 g0592(.A(n655), .B1(n522), .B2(n644), .C1(n533), .C2(n525), .ZN(n656));
  AOI21_X1  g0593(.A(n536), .B1(n656), .B2(n654), .ZN(n657));
  NOR2_X1   g0594(.A1(n657), .A2(n649), .ZN(n658));
  XNOR2_X1  g0595(.A(n658), .B(n648), .ZN(n659));
  AND2_X1   g0596(.A1(375), .A2(103), .ZN(n660));
  XNOR2_X1  g0597(.A(n660), .B(n659), .ZN(n661));
  NOR2_X1   g0598(.A1(n547), .A2(n537), .ZN(n662));
  OAI22_X1  g0599(.A1(n541), .A2(n542), .B1(n435), .B2(n427), .ZN(n663));
  INV_X1    g0600(.A(n536), .ZN(n664));
  AOI21_X1  g0601(.A(n664), .B1(n656), .B2(n654), .ZN(n665));
  AND3_X1   g0602(.A1(n664), .A2(n656), .A3(n654), .ZN(n666));
  OAI221_X1 g0603(.A(n663), .B1(n438), .B2(n437), .C1(n666), .C2(n665), .ZN(n667));
  NAND3_X1  g0604(.A1(n664), .A2(n656), .A3(n654), .ZN(n668));
  OAI221_X1 g0605(.A(n668), .B1(n535), .B2(n657), .C1(n546), .C2(n538), .ZN(n669));
  AOI21_X1  g0606(.A(n549), .B1(n669), .B2(n667), .ZN(n670));
  NOR2_X1   g0607(.A1(n670), .A2(n662), .ZN(n671));
  XNOR2_X1  g0608(.A(n671), .B(n661), .ZN(n672));
  AND2_X1   g0609(.A1(392), .A2(86), .ZN(n673));
  XNOR2_X1  g0610(.A(n673), .B(n672), .ZN(n674));
  NOR2_X1   g0611(.A1(n560), .A2(n550), .ZN(n675));
  OAI22_X1  g0612(.A1(n554), .A2(n555), .B1(n448), .B2(n440), .ZN(n676));
  INV_X1    g0613(.A(n549), .ZN(n677));
  AOI21_X1  g0614(.A(n677), .B1(n669), .B2(n667), .ZN(n678));
  AND3_X1   g0615(.A1(n677), .A2(n669), .A3(n667), .ZN(n679));
  OAI221_X1 g0616(.A(n676), .B1(n451), .B2(n450), .C1(n679), .C2(n678), .ZN(n680));
  NAND3_X1  g0617(.A1(n677), .A2(n669), .A3(n667), .ZN(n681));
  OAI221_X1 g0618(.A(n681), .B1(n548), .B2(n670), .C1(n559), .C2(n551), .ZN(n682));
  AOI21_X1  g0619(.A(n562), .B1(n682), .B2(n680), .ZN(n683));
  NOR2_X1   g0620(.A1(n683), .A2(n675), .ZN(n684));
  XNOR2_X1  g0621(.A(n684), .B(n674), .ZN(n685));
  AND2_X1   g0622(.A1(409), .A2(69), .ZN(n686));
  XNOR2_X1  g0623(.A(n686), .B(n685), .ZN(n687));
  NOR2_X1   g0624(.A1(n573), .A2(n563), .ZN(n688));
  OAI22_X1  g0625(.A1(n567), .A2(n568), .B1(n461), .B2(n453), .ZN(n689));
  INV_X1    g0626(.A(n562), .ZN(n690));
  AOI21_X1  g0627(.A(n690), .B1(n682), .B2(n680), .ZN(n691));
  AND3_X1   g0628(.A1(n690), .A2(n682), .A3(n680), .ZN(n692));
  OAI221_X1 g0629(.A(n689), .B1(n464), .B2(n463), .C1(n692), .C2(n691), .ZN(n693));
  NAND3_X1  g0630(.A1(n690), .A2(n682), .A3(n680), .ZN(n694));
  OAI221_X1 g0631(.A(n694), .B1(n561), .B2(n683), .C1(n572), .C2(n564), .ZN(n695));
  AOI21_X1  g0632(.A(n575), .B1(n695), .B2(n693), .ZN(n696));
  NOR2_X1   g0633(.A1(n696), .A2(n688), .ZN(n697));
  XNOR2_X1  g0634(.A(n697), .B(n687), .ZN(n698));
  AND2_X1   g0635(.A1(426), .A2(52), .ZN(n699));
  XNOR2_X1  g0636(.A(n699), .B(n698), .ZN(n700));
  NOR2_X1   g0637(.A1(n586), .A2(n576), .ZN(n701));
  OAI22_X1  g0638(.A1(n580), .A2(n581), .B1(n474), .B2(n466), .ZN(n702));
  INV_X1    g0639(.A(n575), .ZN(n703));
  AOI21_X1  g0640(.A(n703), .B1(n695), .B2(n693), .ZN(n704));
  AND3_X1   g0641(.A1(n703), .A2(n695), .A3(n693), .ZN(n705));
  OAI221_X1 g0642(.A(n702), .B1(n477), .B2(n476), .C1(n705), .C2(n704), .ZN(n706));
  NAND3_X1  g0643(.A1(n703), .A2(n695), .A3(n693), .ZN(n707));
  OAI221_X1 g0644(.A(n707), .B1(n574), .B2(n696), .C1(n585), .C2(n577), .ZN(n708));
  AOI21_X1  g0645(.A(n588), .B1(n708), .B2(n706), .ZN(n709));
  NOR2_X1   g0646(.A1(n709), .A2(n701), .ZN(n710));
  XNOR2_X1  g0647(.A(n710), .B(n700), .ZN(n711));
  AND2_X1   g0648(.A1(443), .A2(35), .ZN(n712));
  XNOR2_X1  g0649(.A(n712), .B(n711), .ZN(n713));
  NOR2_X1   g0650(.A1(n599), .A2(n589), .ZN(n714));
  OAI22_X1  g0651(.A1(n593), .A2(n594), .B1(n487), .B2(n479), .ZN(n715));
  INV_X1    g0652(.A(n588), .ZN(n716));
  AOI21_X1  g0653(.A(n716), .B1(n708), .B2(n706), .ZN(n717));
  AND3_X1   g0654(.A1(n716), .A2(n708), .A3(n706), .ZN(n718));
  OAI221_X1 g0655(.A(n715), .B1(n490), .B2(n489), .C1(n718), .C2(n717), .ZN(n719));
  NAND3_X1  g0656(.A1(n716), .A2(n708), .A3(n706), .ZN(n720));
  OAI221_X1 g0657(.A(n720), .B1(n587), .B2(n709), .C1(n598), .C2(n590), .ZN(n721));
  AOI21_X1  g0658(.A(n601), .B1(n721), .B2(n719), .ZN(n722));
  NOR2_X1   g0659(.A1(n722), .A2(n714), .ZN(n723));
  XNOR2_X1  g0660(.A(n723), .B(n713), .ZN(n724));
  AND2_X1   g0661(.A1(460), .A2(18), .ZN(n725));
  XNOR2_X1  g0662(.A(n725), .B(n724), .ZN(n726));
  NOR2_X1   g0663(.A1(n604), .A2(n602), .ZN(n727));
  AOI21_X1  g0664(.A(n727), .B1(n607), .B2(n605), .ZN(n728));
  XOR2_X1   g0665(.A(n728), .B(n726), .ZN(n729));
  AND2_X1   g0666(.A1(477), .A2(\1 ), .ZN(n730));
  INV_X1    g0667(.A(n730), .ZN(n731));
  XNOR2_X1  g0668(.A(n731), .B(n729), .ZN(5308));
  AND4_X1   g0669(.A1(273), .A2(222), .A3(205), .A4(290), .ZN(n733));
  AOI22_X1  g0670(.A1(273), .A2(222), .B1(205), .B2(290), .ZN(n734));
  NOR2_X1   g0671(.A1(n734), .A2(n733), .ZN(n735));
  XNOR2_X1  g0672(.A(n735), .B(n609), .ZN(n736));
  AND2_X1   g0673(.A1(307), .A2(188), .ZN(n737));
  XNOR2_X1  g0674(.A(n737), .B(n736), .ZN(n738));
  NOR2_X1   g0675(.A1(n611), .A2(n498), .ZN(n739));
  OAI21_X1  g0676(.A(n498), .B1(n610), .B2(n609), .ZN(n740));
  OR3_X1    g0677(.A1(n610), .A2(n609), .A3(n498), .ZN(n741));
  AOI21_X1  g0678(.A(n613), .B1(n741), .B2(n740), .ZN(n742));
  NOR2_X1   g0679(.A1(n742), .A2(n739), .ZN(n743));
  XNOR2_X1  g0680(.A(n743), .B(n738), .ZN(n744));
  AND2_X1   g0681(.A1(324), .A2(171), .ZN(n745));
  XNOR2_X1  g0682(.A(n745), .B(n744), .ZN(n746));
  NOR2_X1   g0683(.A1(n619), .A2(n614), .ZN(n747));
  OR2_X1    g0684(.A1(n500), .A2(n400), .ZN(n748));
  NAND2_X1  g0685(.A1(307), .A2(171), .ZN(n749));
  AOI21_X1  g0686(.A(n749), .B1(n741), .B2(n740), .ZN(n750));
  AND3_X1   g0687(.A1(n749), .A2(n741), .A3(n740), .ZN(n751));
  OAI221_X1 g0688(.A(n748), .B1(n502), .B2(n501), .C1(n751), .C2(n750), .ZN(n752));
  NAND3_X1  g0689(.A1(n749), .A2(n741), .A3(n740), .ZN(n753));
  OAI221_X1 g0690(.A(n753), .B1(n612), .B2(n742), .C1(n618), .C2(n615), .ZN(n754));
  AOI21_X1  g0691(.A(n621), .B1(n754), .B2(n752), .ZN(n755));
  NOR2_X1   g0692(.A1(n755), .A2(n747), .ZN(n756));
  XNOR2_X1  g0693(.A(n756), .B(n746), .ZN(n757));
  AND2_X1   g0694(.A1(341), .A2(154), .ZN(n758));
  XNOR2_X1  g0695(.A(n758), .B(n757), .ZN(n759));
  NOR2_X1   g0696(.A1(n632), .A2(n622), .ZN(n760));
  OAI22_X1  g0697(.A1(n626), .A2(n627), .B1(n507), .B2(n504), .ZN(n761));
  INV_X1    g0698(.A(n621), .ZN(n762));
  AOI21_X1  g0699(.A(n762), .B1(n754), .B2(n752), .ZN(n763));
  AND3_X1   g0700(.A1(n762), .A2(n754), .A3(n752), .ZN(n764));
  OAI221_X1 g0701(.A(n761), .B1(n510), .B2(n509), .C1(n764), .C2(n763), .ZN(n765));
  NAND3_X1  g0702(.A1(n762), .A2(n754), .A3(n752), .ZN(n766));
  OAI221_X1 g0703(.A(n766), .B1(n620), .B2(n755), .C1(n631), .C2(n623), .ZN(n767));
  AOI21_X1  g0704(.A(n634), .B1(n767), .B2(n765), .ZN(n768));
  NOR2_X1   g0705(.A1(n768), .A2(n760), .ZN(n769));
  XNOR2_X1  g0706(.A(n769), .B(n759), .ZN(n770));
  AND2_X1   g0707(.A1(358), .A2(137), .ZN(n771));
  XNOR2_X1  g0708(.A(n771), .B(n770), .ZN(n772));
  NOR2_X1   g0709(.A1(n645), .A2(n635), .ZN(n773));
  OAI22_X1  g0710(.A1(n639), .A2(n640), .B1(n520), .B2(n512), .ZN(n774));
  INV_X1    g0711(.A(n634), .ZN(n775));
  AOI21_X1  g0712(.A(n775), .B1(n767), .B2(n765), .ZN(n776));
  AND3_X1   g0713(.A1(n775), .A2(n767), .A3(n765), .ZN(n777));
  OAI221_X1 g0714(.A(n774), .B1(n523), .B2(n522), .C1(n777), .C2(n776), .ZN(n778));
  NAND3_X1  g0715(.A1(n775), .A2(n767), .A3(n765), .ZN(n779));
  OAI221_X1 g0716(.A(n779), .B1(n633), .B2(n768), .C1(n644), .C2(n636), .ZN(n780));
  AOI21_X1  g0717(.A(n647), .B1(n780), .B2(n778), .ZN(n781));
  NOR2_X1   g0718(.A1(n781), .A2(n773), .ZN(n782));
  XNOR2_X1  g0719(.A(n782), .B(n772), .ZN(n783));
  AND2_X1   g0720(.A1(375), .A2(120), .ZN(n784));
  XNOR2_X1  g0721(.A(n784), .B(n783), .ZN(n785));
  NOR2_X1   g0722(.A1(n658), .A2(n648), .ZN(n786));
  OAI22_X1  g0723(.A1(n652), .A2(n653), .B1(n533), .B2(n525), .ZN(n787));
  INV_X1    g0724(.A(n647), .ZN(n788));
  AOI21_X1  g0725(.A(n788), .B1(n780), .B2(n778), .ZN(n789));
  AND3_X1   g0726(.A1(n788), .A2(n780), .A3(n778), .ZN(n790));
  OAI221_X1 g0727(.A(n787), .B1(n536), .B2(n535), .C1(n790), .C2(n789), .ZN(n791));
  NAND3_X1  g0728(.A1(n788), .A2(n780), .A3(n778), .ZN(n792));
  OAI221_X1 g0729(.A(n792), .B1(n646), .B2(n781), .C1(n657), .C2(n649), .ZN(n793));
  AOI21_X1  g0730(.A(n660), .B1(n793), .B2(n791), .ZN(n794));
  NOR2_X1   g0731(.A1(n794), .A2(n786), .ZN(n795));
  XNOR2_X1  g0732(.A(n795), .B(n785), .ZN(n796));
  AND2_X1   g0733(.A1(392), .A2(103), .ZN(n797));
  XNOR2_X1  g0734(.A(n797), .B(n796), .ZN(n798));
  NOR2_X1   g0735(.A1(n671), .A2(n661), .ZN(n799));
  OAI22_X1  g0736(.A1(n665), .A2(n666), .B1(n546), .B2(n538), .ZN(n800));
  INV_X1    g0737(.A(n660), .ZN(n801));
  AOI21_X1  g0738(.A(n801), .B1(n793), .B2(n791), .ZN(n802));
  AND3_X1   g0739(.A1(n801), .A2(n793), .A3(n791), .ZN(n803));
  OAI221_X1 g0740(.A(n800), .B1(n549), .B2(n548), .C1(n803), .C2(n802), .ZN(n804));
  NAND3_X1  g0741(.A1(n801), .A2(n793), .A3(n791), .ZN(n805));
  OAI221_X1 g0742(.A(n805), .B1(n659), .B2(n794), .C1(n670), .C2(n662), .ZN(n806));
  AOI21_X1  g0743(.A(n673), .B1(n806), .B2(n804), .ZN(n807));
  NOR2_X1   g0744(.A1(n807), .A2(n799), .ZN(n808));
  XNOR2_X1  g0745(.A(n808), .B(n798), .ZN(n809));
  AND2_X1   g0746(.A1(409), .A2(86), .ZN(n810));
  XNOR2_X1  g0747(.A(n810), .B(n809), .ZN(n811));
  NOR2_X1   g0748(.A1(n684), .A2(n674), .ZN(n812));
  OAI22_X1  g0749(.A1(n678), .A2(n679), .B1(n559), .B2(n551), .ZN(n813));
  INV_X1    g0750(.A(n673), .ZN(n814));
  AOI21_X1  g0751(.A(n814), .B1(n806), .B2(n804), .ZN(n815));
  AND3_X1   g0752(.A1(n814), .A2(n806), .A3(n804), .ZN(n816));
  OAI221_X1 g0753(.A(n813), .B1(n562), .B2(n561), .C1(n816), .C2(n815), .ZN(n817));
  NAND3_X1  g0754(.A1(n814), .A2(n806), .A3(n804), .ZN(n818));
  OAI221_X1 g0755(.A(n818), .B1(n672), .B2(n807), .C1(n683), .C2(n675), .ZN(n819));
  AOI21_X1  g0756(.A(n686), .B1(n819), .B2(n817), .ZN(n820));
  NOR2_X1   g0757(.A1(n820), .A2(n812), .ZN(n821));
  XNOR2_X1  g0758(.A(n821), .B(n811), .ZN(n822));
  AND2_X1   g0759(.A1(426), .A2(69), .ZN(n823));
  XNOR2_X1  g0760(.A(n823), .B(n822), .ZN(n824));
  NOR2_X1   g0761(.A1(n697), .A2(n687), .ZN(n825));
  OAI22_X1  g0762(.A1(n691), .A2(n692), .B1(n572), .B2(n564), .ZN(n826));
  INV_X1    g0763(.A(n686), .ZN(n827));
  AOI21_X1  g0764(.A(n827), .B1(n819), .B2(n817), .ZN(n828));
  AND3_X1   g0765(.A1(n827), .A2(n819), .A3(n817), .ZN(n829));
  OAI221_X1 g0766(.A(n826), .B1(n575), .B2(n574), .C1(n829), .C2(n828), .ZN(n830));
  NAND3_X1  g0767(.A1(n827), .A2(n819), .A3(n817), .ZN(n831));
  OAI221_X1 g0768(.A(n831), .B1(n685), .B2(n820), .C1(n696), .C2(n688), .ZN(n832));
  AOI21_X1  g0769(.A(n699), .B1(n832), .B2(n830), .ZN(n833));
  NOR2_X1   g0770(.A1(n833), .A2(n825), .ZN(n834));
  XNOR2_X1  g0771(.A(n834), .B(n824), .ZN(n835));
  AND2_X1   g0772(.A1(443), .A2(52), .ZN(n836));
  XNOR2_X1  g0773(.A(n836), .B(n835), .ZN(n837));
  NOR2_X1   g0774(.A1(n710), .A2(n700), .ZN(n838));
  OAI22_X1  g0775(.A1(n704), .A2(n705), .B1(n585), .B2(n577), .ZN(n839));
  INV_X1    g0776(.A(n699), .ZN(n840));
  AOI21_X1  g0777(.A(n840), .B1(n832), .B2(n830), .ZN(n841));
  AND3_X1   g0778(.A1(n840), .A2(n832), .A3(n830), .ZN(n842));
  OAI221_X1 g0779(.A(n839), .B1(n588), .B2(n587), .C1(n842), .C2(n841), .ZN(n843));
  NAND3_X1  g0780(.A1(n840), .A2(n832), .A3(n830), .ZN(n844));
  OAI221_X1 g0781(.A(n844), .B1(n698), .B2(n833), .C1(n709), .C2(n701), .ZN(n845));
  AOI21_X1  g0782(.A(n712), .B1(n845), .B2(n843), .ZN(n846));
  NOR2_X1   g0783(.A1(n846), .A2(n838), .ZN(n847));
  XNOR2_X1  g0784(.A(n847), .B(n837), .ZN(n848));
  AND2_X1   g0785(.A1(460), .A2(35), .ZN(n849));
  XNOR2_X1  g0786(.A(n849), .B(n848), .ZN(n850));
  NOR2_X1   g0787(.A1(n723), .A2(n713), .ZN(n851));
  OAI22_X1  g0788(.A1(n717), .A2(n718), .B1(n598), .B2(n590), .ZN(n852));
  INV_X1    g0789(.A(n712), .ZN(n853));
  AOI21_X1  g0790(.A(n853), .B1(n845), .B2(n843), .ZN(n854));
  AND3_X1   g0791(.A1(n853), .A2(n845), .A3(n843), .ZN(n855));
  OAI221_X1 g0792(.A(n852), .B1(n601), .B2(n600), .C1(n855), .C2(n854), .ZN(n856));
  NAND3_X1  g0793(.A1(n853), .A2(n845), .A3(n843), .ZN(n857));
  OAI221_X1 g0794(.A(n857), .B1(n711), .B2(n846), .C1(n722), .C2(n714), .ZN(n858));
  AOI21_X1  g0795(.A(n725), .B1(n858), .B2(n856), .ZN(n859));
  NOR2_X1   g0796(.A1(n859), .A2(n851), .ZN(n860));
  XNOR2_X1  g0797(.A(n860), .B(n850), .ZN(n861));
  AND2_X1   g0798(.A1(477), .A2(18), .ZN(n862));
  XNOR2_X1  g0799(.A(n862), .B(n861), .ZN(n863));
  NOR2_X1   g0800(.A1(n728), .A2(n726), .ZN(n864));
  AOI21_X1  g0801(.A(n864), .B1(n731), .B2(n729), .ZN(n865));
  XOR2_X1   g0802(.A(n865), .B(n863), .ZN(n866));
  AND2_X1   g0803(.A1(494), .A2(\1 ), .ZN(n867));
  INV_X1    g0804(.A(n867), .ZN(n868));
  XNOR2_X1  g0805(.A(n868), .B(n866), .ZN(5672));
  AND4_X1   g0806(.A1(273), .A2(239), .A3(222), .A4(290), .ZN(n870));
  AOI22_X1  g0807(.A1(273), .A2(239), .B1(222), .B2(290), .ZN(n871));
  NOR2_X1   g0808(.A1(n871), .A2(n870), .ZN(n872));
  XNOR2_X1  g0809(.A(n872), .B(n733), .ZN(n873));
  AND2_X1   g0810(.A1(307), .A2(205), .ZN(n874));
  XNOR2_X1  g0811(.A(n874), .B(n873), .ZN(n875));
  NOR2_X1   g0812(.A1(n735), .A2(n609), .ZN(n876));
  OAI21_X1  g0813(.A(n609), .B1(n734), .B2(n733), .ZN(n877));
  OR3_X1    g0814(.A1(n734), .A2(n733), .A3(n609), .ZN(n878));
  AOI21_X1  g0815(.A(n737), .B1(n878), .B2(n877), .ZN(n879));
  NOR2_X1   g0816(.A1(n879), .A2(n876), .ZN(n880));
  XNOR2_X1  g0817(.A(n880), .B(n875), .ZN(n881));
  AND2_X1   g0818(.A1(324), .A2(188), .ZN(n882));
  XNOR2_X1  g0819(.A(n882), .B(n881), .ZN(n883));
  NOR2_X1   g0820(.A1(n743), .A2(n738), .ZN(n884));
  OR2_X1    g0821(.A1(n611), .A2(n498), .ZN(n885));
  NAND2_X1  g0822(.A1(307), .A2(188), .ZN(n886));
  AOI21_X1  g0823(.A(n886), .B1(n878), .B2(n877), .ZN(n887));
  AND3_X1   g0824(.A1(n886), .A2(n878), .A3(n877), .ZN(n888));
  OAI221_X1 g0825(.A(n885), .B1(n613), .B2(n612), .C1(n888), .C2(n887), .ZN(n889));
  NAND3_X1  g0826(.A1(n886), .A2(n878), .A3(n877), .ZN(n890));
  OAI221_X1 g0827(.A(n890), .B1(n736), .B2(n879), .C1(n742), .C2(n739), .ZN(n891));
  AOI21_X1  g0828(.A(n745), .B1(n891), .B2(n889), .ZN(n892));
  NOR2_X1   g0829(.A1(n892), .A2(n884), .ZN(n893));
  XNOR2_X1  g0830(.A(n893), .B(n883), .ZN(n894));
  AND2_X1   g0831(.A1(341), .A2(171), .ZN(n895));
  XNOR2_X1  g0832(.A(n895), .B(n894), .ZN(n896));
  NOR2_X1   g0833(.A1(n756), .A2(n746), .ZN(n897));
  OAI22_X1  g0834(.A1(n750), .A2(n751), .B1(n618), .B2(n615), .ZN(n898));
  INV_X1    g0835(.A(n745), .ZN(n899));
  AOI21_X1  g0836(.A(n899), .B1(n891), .B2(n889), .ZN(n900));
  AND3_X1   g0837(.A1(n899), .A2(n891), .A3(n889), .ZN(n901));
  OAI221_X1 g0838(.A(n898), .B1(n621), .B2(n620), .C1(n901), .C2(n900), .ZN(n902));
  NAND3_X1  g0839(.A1(n899), .A2(n891), .A3(n889), .ZN(n903));
  OAI221_X1 g0840(.A(n903), .B1(n744), .B2(n892), .C1(n755), .C2(n747), .ZN(n904));
  AOI21_X1  g0841(.A(n758), .B1(n904), .B2(n902), .ZN(n905));
  NOR2_X1   g0842(.A1(n905), .A2(n897), .ZN(n906));
  XNOR2_X1  g0843(.A(n906), .B(n896), .ZN(n907));
  AND2_X1   g0844(.A1(358), .A2(154), .ZN(n908));
  XNOR2_X1  g0845(.A(n908), .B(n907), .ZN(n909));
  NOR2_X1   g0846(.A1(n769), .A2(n759), .ZN(n910));
  OAI22_X1  g0847(.A1(n763), .A2(n764), .B1(n631), .B2(n623), .ZN(n911));
  INV_X1    g0848(.A(n758), .ZN(n912));
  AOI21_X1  g0849(.A(n912), .B1(n904), .B2(n902), .ZN(n913));
  AND3_X1   g0850(.A1(n912), .A2(n904), .A3(n902), .ZN(n914));
  OAI221_X1 g0851(.A(n911), .B1(n634), .B2(n633), .C1(n914), .C2(n913), .ZN(n915));
  NAND3_X1  g0852(.A1(n912), .A2(n904), .A3(n902), .ZN(n916));
  OAI221_X1 g0853(.A(n916), .B1(n757), .B2(n905), .C1(n768), .C2(n760), .ZN(n917));
  AOI21_X1  g0854(.A(n771), .B1(n917), .B2(n915), .ZN(n918));
  NOR2_X1   g0855(.A1(n918), .A2(n910), .ZN(n919));
  XNOR2_X1  g0856(.A(n919), .B(n909), .ZN(n920));
  AND2_X1   g0857(.A1(375), .A2(137), .ZN(n921));
  XNOR2_X1  g0858(.A(n921), .B(n920), .ZN(n922));
  NOR2_X1   g0859(.A1(n782), .A2(n772), .ZN(n923));
  OAI22_X1  g0860(.A1(n776), .A2(n777), .B1(n644), .B2(n636), .ZN(n924));
  INV_X1    g0861(.A(n771), .ZN(n925));
  AOI21_X1  g0862(.A(n925), .B1(n917), .B2(n915), .ZN(n926));
  AND3_X1   g0863(.A1(n925), .A2(n917), .A3(n915), .ZN(n927));
  OAI221_X1 g0864(.A(n924), .B1(n647), .B2(n646), .C1(n927), .C2(n926), .ZN(n928));
  NAND3_X1  g0865(.A1(n925), .A2(n917), .A3(n915), .ZN(n929));
  OAI221_X1 g0866(.A(n929), .B1(n770), .B2(n918), .C1(n781), .C2(n773), .ZN(n930));
  AOI21_X1  g0867(.A(n784), .B1(n930), .B2(n928), .ZN(n931));
  NOR2_X1   g0868(.A1(n931), .A2(n923), .ZN(n932));
  XNOR2_X1  g0869(.A(n932), .B(n922), .ZN(n933));
  AND2_X1   g0870(.A1(392), .A2(120), .ZN(n934));
  XNOR2_X1  g0871(.A(n934), .B(n933), .ZN(n935));
  NOR2_X1   g0872(.A1(n795), .A2(n785), .ZN(n936));
  OAI22_X1  g0873(.A1(n789), .A2(n790), .B1(n657), .B2(n649), .ZN(n937));
  INV_X1    g0874(.A(n784), .ZN(n938));
  AOI21_X1  g0875(.A(n938), .B1(n930), .B2(n928), .ZN(n939));
  AND3_X1   g0876(.A1(n938), .A2(n930), .A3(n928), .ZN(n940));
  OAI221_X1 g0877(.A(n937), .B1(n660), .B2(n659), .C1(n940), .C2(n939), .ZN(n941));
  NAND3_X1  g0878(.A1(n938), .A2(n930), .A3(n928), .ZN(n942));
  OAI221_X1 g0879(.A(n942), .B1(n783), .B2(n931), .C1(n794), .C2(n786), .ZN(n943));
  AOI21_X1  g0880(.A(n797), .B1(n943), .B2(n941), .ZN(n944));
  NOR2_X1   g0881(.A1(n944), .A2(n936), .ZN(n945));
  XNOR2_X1  g0882(.A(n945), .B(n935), .ZN(n946));
  AND2_X1   g0883(.A1(409), .A2(103), .ZN(n947));
  XNOR2_X1  g0884(.A(n947), .B(n946), .ZN(n948));
  NOR2_X1   g0885(.A1(n808), .A2(n798), .ZN(n949));
  OAI22_X1  g0886(.A1(n802), .A2(n803), .B1(n670), .B2(n662), .ZN(n950));
  INV_X1    g0887(.A(n797), .ZN(n951));
  AOI21_X1  g0888(.A(n951), .B1(n943), .B2(n941), .ZN(n952));
  AND3_X1   g0889(.A1(n951), .A2(n943), .A3(n941), .ZN(n953));
  OAI221_X1 g0890(.A(n950), .B1(n673), .B2(n672), .C1(n953), .C2(n952), .ZN(n954));
  NAND3_X1  g0891(.A1(n951), .A2(n943), .A3(n941), .ZN(n955));
  OAI221_X1 g0892(.A(n955), .B1(n796), .B2(n944), .C1(n807), .C2(n799), .ZN(n956));
  AOI21_X1  g0893(.A(n810), .B1(n956), .B2(n954), .ZN(n957));
  NOR2_X1   g0894(.A1(n957), .A2(n949), .ZN(n958));
  XNOR2_X1  g0895(.A(n958), .B(n948), .ZN(n959));
  AND2_X1   g0896(.A1(426), .A2(86), .ZN(n960));
  XNOR2_X1  g0897(.A(n960), .B(n959), .ZN(n961));
  NOR2_X1   g0898(.A1(n821), .A2(n811), .ZN(n962));
  OAI22_X1  g0899(.A1(n815), .A2(n816), .B1(n683), .B2(n675), .ZN(n963));
  INV_X1    g0900(.A(n810), .ZN(n964));
  AOI21_X1  g0901(.A(n964), .B1(n956), .B2(n954), .ZN(n965));
  AND3_X1   g0902(.A1(n964), .A2(n956), .A3(n954), .ZN(n966));
  OAI221_X1 g0903(.A(n963), .B1(n686), .B2(n685), .C1(n966), .C2(n965), .ZN(n967));
  NAND3_X1  g0904(.A1(n964), .A2(n956), .A3(n954), .ZN(n968));
  OAI221_X1 g0905(.A(n968), .B1(n809), .B2(n957), .C1(n820), .C2(n812), .ZN(n969));
  AOI21_X1  g0906(.A(n823), .B1(n969), .B2(n967), .ZN(n970));
  NOR2_X1   g0907(.A1(n970), .A2(n962), .ZN(n971));
  XNOR2_X1  g0908(.A(n971), .B(n961), .ZN(n972));
  AND2_X1   g0909(.A1(443), .A2(69), .ZN(n973));
  XNOR2_X1  g0910(.A(n973), .B(n972), .ZN(n974));
  NOR2_X1   g0911(.A1(n834), .A2(n824), .ZN(n975));
  OAI22_X1  g0912(.A1(n828), .A2(n829), .B1(n696), .B2(n688), .ZN(n976));
  INV_X1    g0913(.A(n823), .ZN(n977));
  AOI21_X1  g0914(.A(n977), .B1(n969), .B2(n967), .ZN(n978));
  AND3_X1   g0915(.A1(n977), .A2(n969), .A3(n967), .ZN(n979));
  OAI221_X1 g0916(.A(n976), .B1(n699), .B2(n698), .C1(n979), .C2(n978), .ZN(n980));
  NAND3_X1  g0917(.A1(n977), .A2(n969), .A3(n967), .ZN(n981));
  OAI221_X1 g0918(.A(n981), .B1(n822), .B2(n970), .C1(n833), .C2(n825), .ZN(n982));
  AOI21_X1  g0919(.A(n836), .B1(n982), .B2(n980), .ZN(n983));
  NOR2_X1   g0920(.A1(n983), .A2(n975), .ZN(n984));
  XNOR2_X1  g0921(.A(n984), .B(n974), .ZN(n985));
  AND2_X1   g0922(.A1(460), .A2(52), .ZN(n986));
  XNOR2_X1  g0923(.A(n986), .B(n985), .ZN(n987));
  NOR2_X1   g0924(.A1(n847), .A2(n837), .ZN(n988));
  OAI22_X1  g0925(.A1(n841), .A2(n842), .B1(n709), .B2(n701), .ZN(n989));
  INV_X1    g0926(.A(n836), .ZN(n990));
  AOI21_X1  g0927(.A(n990), .B1(n982), .B2(n980), .ZN(n991));
  AND3_X1   g0928(.A1(n990), .A2(n982), .A3(n980), .ZN(n992));
  OAI221_X1 g0929(.A(n989), .B1(n712), .B2(n711), .C1(n992), .C2(n991), .ZN(n993));
  NAND3_X1  g0930(.A1(n990), .A2(n982), .A3(n980), .ZN(n994));
  OAI221_X1 g0931(.A(n994), .B1(n835), .B2(n983), .C1(n846), .C2(n838), .ZN(n995));
  AOI21_X1  g0932(.A(n849), .B1(n995), .B2(n993), .ZN(n996));
  NOR2_X1   g0933(.A1(n996), .A2(n988), .ZN(n997));
  XNOR2_X1  g0934(.A(n997), .B(n987), .ZN(n998));
  AND2_X1   g0935(.A1(477), .A2(35), .ZN(n999));
  XNOR2_X1  g0936(.A(n999), .B(n998), .ZN(n1000));
  NOR2_X1   g0937(.A1(n860), .A2(n850), .ZN(n1001));
  OAI22_X1  g0938(.A1(n854), .A2(n855), .B1(n722), .B2(n714), .ZN(n1002));
  INV_X1    g0939(.A(n849), .ZN(n1003));
  AOI21_X1  g0940(.A(n1003), .B1(n995), .B2(n993), .ZN(n1004));
  AND3_X1   g0941(.A1(n1003), .A2(n995), .A3(n993), .ZN(n1005));
  OAI221_X1 g0942(.A(n1002), .B1(n725), .B2(n724), .C1(n1005), .C2(n1004), .ZN(n1006));
  NAND3_X1  g0943(.A1(n1003), .A2(n995), .A3(n993), .ZN(n1007));
  OAI221_X1 g0944(.A(n1007), .B1(n848), .B2(n996), .C1(n859), .C2(n851), .ZN(n1008));
  AOI21_X1  g0945(.A(n862), .B1(n1008), .B2(n1006), .ZN(n1009));
  NOR2_X1   g0946(.A1(n1009), .A2(n1001), .ZN(n1010));
  XNOR2_X1  g0947(.A(n1010), .B(n1000), .ZN(n1011));
  AND2_X1   g0948(.A1(494), .A2(18), .ZN(n1012));
  XNOR2_X1  g0949(.A(n1012), .B(n1011), .ZN(n1013));
  NOR2_X1   g0950(.A1(n865), .A2(n863), .ZN(n1014));
  AOI21_X1  g0951(.A(n1014), .B1(n868), .B2(n866), .ZN(n1015));
  XOR2_X1   g0952(.A(n1015), .B(n1013), .ZN(n1016));
  AND2_X1   g0953(.A1(511), .A2(\1 ), .ZN(n1017));
  INV_X1    g0954(.A(n1017), .ZN(n1018));
  XNOR2_X1  g0955(.A(n1018), .B(n1016), .ZN(5971));
  AND4_X1   g0956(.A1(273), .A2(256), .A3(239), .A4(290), .ZN(n1020));
  AOI22_X1  g0957(.A1(273), .A2(256), .B1(239), .B2(290), .ZN(n1021));
  NOR2_X1   g0958(.A1(n1021), .A2(n1020), .ZN(n1022));
  XNOR2_X1  g0959(.A(n1022), .B(n870), .ZN(n1023));
  AND2_X1   g0960(.A1(307), .A2(222), .ZN(n1024));
  XNOR2_X1  g0961(.A(n1024), .B(n1023), .ZN(n1025));
  NOR2_X1   g0962(.A1(n872), .A2(n733), .ZN(n1026));
  OAI21_X1  g0963(.A(n733), .B1(n871), .B2(n870), .ZN(n1027));
  OR3_X1    g0964(.A1(n871), .A2(n870), .A3(n733), .ZN(n1028));
  AOI21_X1  g0965(.A(n874), .B1(n1028), .B2(n1027), .ZN(n1029));
  NOR2_X1   g0966(.A1(n1029), .A2(n1026), .ZN(n1030));
  XNOR2_X1  g0967(.A(n1030), .B(n1025), .ZN(n1031));
  AND2_X1   g0968(.A1(324), .A2(205), .ZN(n1032));
  XNOR2_X1  g0969(.A(n1032), .B(n1031), .ZN(n1033));
  NOR2_X1   g0970(.A1(n880), .A2(n875), .ZN(n1034));
  OR2_X1    g0971(.A1(n735), .A2(n609), .ZN(n1035));
  NAND2_X1  g0972(.A1(307), .A2(205), .ZN(n1036));
  AOI21_X1  g0973(.A(n1036), .B1(n1028), .B2(n1027), .ZN(n1037));
  AND3_X1   g0974(.A1(n1036), .A2(n1028), .A3(n1027), .ZN(n1038));
  OAI221_X1 g0975(.A(n1035), .B1(n737), .B2(n736), .C1(n1038), .C2(n1037), .ZN(n1039));
  NAND3_X1  g0976(.A1(n1036), .A2(n1028), .A3(n1027), .ZN(n1040));
  OAI221_X1 g0977(.A(n1040), .B1(n873), .B2(n1029), .C1(n879), .C2(n876), .ZN(n1041));
  AOI21_X1  g0978(.A(n882), .B1(n1041), .B2(n1039), .ZN(n1042));
  NOR2_X1   g0979(.A1(n1042), .A2(n1034), .ZN(n1043));
  XNOR2_X1  g0980(.A(n1043), .B(n1033), .ZN(n1044));
  AND2_X1   g0981(.A1(341), .A2(188), .ZN(n1045));
  XNOR2_X1  g0982(.A(n1045), .B(n1044), .ZN(n1046));
  NOR2_X1   g0983(.A1(n893), .A2(n883), .ZN(n1047));
  OAI22_X1  g0984(.A1(n887), .A2(n888), .B1(n742), .B2(n739), .ZN(n1048));
  INV_X1    g0985(.A(n882), .ZN(n1049));
  AOI21_X1  g0986(.A(n1049), .B1(n1041), .B2(n1039), .ZN(n1050));
  AND3_X1   g0987(.A1(n1049), .A2(n1041), .A3(n1039), .ZN(n1051));
  OAI221_X1 g0988(.A(n1048), .B1(n745), .B2(n744), .C1(n1051), .C2(n1050), .ZN(n1052));
  NAND3_X1  g0989(.A1(n1049), .A2(n1041), .A3(n1039), .ZN(n1053));
  OAI221_X1 g0990(.A(n1053), .B1(n881), .B2(n1042), .C1(n892), .C2(n884), .ZN(n1054));
  AOI21_X1  g0991(.A(n895), .B1(n1054), .B2(n1052), .ZN(n1055));
  NOR2_X1   g0992(.A1(n1055), .A2(n1047), .ZN(n1056));
  XNOR2_X1  g0993(.A(n1056), .B(n1046), .ZN(n1057));
  AND2_X1   g0994(.A1(358), .A2(171), .ZN(n1058));
  XNOR2_X1  g0995(.A(n1058), .B(n1057), .ZN(n1059));
  NOR2_X1   g0996(.A1(n906), .A2(n896), .ZN(n1060));
  OAI22_X1  g0997(.A1(n900), .A2(n901), .B1(n755), .B2(n747), .ZN(n1061));
  INV_X1    g0998(.A(n895), .ZN(n1062));
  AOI21_X1  g0999(.A(n1062), .B1(n1054), .B2(n1052), .ZN(n1063));
  AND3_X1   g1000(.A1(n1062), .A2(n1054), .A3(n1052), .ZN(n1064));
  OAI221_X1 g1001(.A(n1061), .B1(n758), .B2(n757), .C1(n1064), .C2(n1063), .ZN(n1065));
  NAND3_X1  g1002(.A1(n1062), .A2(n1054), .A3(n1052), .ZN(n1066));
  OAI221_X1 g1003(.A(n1066), .B1(n894), .B2(n1055), .C1(n905), .C2(n897), .ZN(n1067));
  AOI21_X1  g1004(.A(n908), .B1(n1067), .B2(n1065), .ZN(n1068));
  NOR2_X1   g1005(.A1(n1068), .A2(n1060), .ZN(n1069));
  XNOR2_X1  g1006(.A(n1069), .B(n1059), .ZN(n1070));
  AND2_X1   g1007(.A1(375), .A2(154), .ZN(n1071));
  XNOR2_X1  g1008(.A(n1071), .B(n1070), .ZN(n1072));
  NOR2_X1   g1009(.A1(n919), .A2(n909), .ZN(n1073));
  OAI22_X1  g1010(.A1(n913), .A2(n914), .B1(n768), .B2(n760), .ZN(n1074));
  INV_X1    g1011(.A(n908), .ZN(n1075));
  AOI21_X1  g1012(.A(n1075), .B1(n1067), .B2(n1065), .ZN(n1076));
  AND3_X1   g1013(.A1(n1075), .A2(n1067), .A3(n1065), .ZN(n1077));
  OAI221_X1 g1014(.A(n1074), .B1(n771), .B2(n770), .C1(n1077), .C2(n1076), .ZN(n1078));
  NAND3_X1  g1015(.A1(n1075), .A2(n1067), .A3(n1065), .ZN(n1079));
  OAI221_X1 g1016(.A(n1079), .B1(n907), .B2(n1068), .C1(n918), .C2(n910), .ZN(n1080));
  AOI21_X1  g1017(.A(n921), .B1(n1080), .B2(n1078), .ZN(n1081));
  NOR2_X1   g1018(.A1(n1081), .A2(n1073), .ZN(n1082));
  XNOR2_X1  g1019(.A(n1082), .B(n1072), .ZN(n1083));
  AND2_X1   g1020(.A1(392), .A2(137), .ZN(n1084));
  XNOR2_X1  g1021(.A(n1084), .B(n1083), .ZN(n1085));
  NOR2_X1   g1022(.A1(n932), .A2(n922), .ZN(n1086));
  OAI22_X1  g1023(.A1(n926), .A2(n927), .B1(n781), .B2(n773), .ZN(n1087));
  INV_X1    g1024(.A(n921), .ZN(n1088));
  AOI21_X1  g1025(.A(n1088), .B1(n1080), .B2(n1078), .ZN(n1089));
  AND3_X1   g1026(.A1(n1088), .A2(n1080), .A3(n1078), .ZN(n1090));
  OAI221_X1 g1027(.A(n1087), .B1(n784), .B2(n783), .C1(n1090), .C2(n1089), .ZN(n1091));
  NAND3_X1  g1028(.A1(n1088), .A2(n1080), .A3(n1078), .ZN(n1092));
  OAI221_X1 g1029(.A(n1092), .B1(n920), .B2(n1081), .C1(n931), .C2(n923), .ZN(n1093));
  AOI21_X1  g1030(.A(n934), .B1(n1093), .B2(n1091), .ZN(n1094));
  NOR2_X1   g1031(.A1(n1094), .A2(n1086), .ZN(n1095));
  XNOR2_X1  g1032(.A(n1095), .B(n1085), .ZN(n1096));
  AND2_X1   g1033(.A1(409), .A2(120), .ZN(n1097));
  XNOR2_X1  g1034(.A(n1097), .B(n1096), .ZN(n1098));
  NOR2_X1   g1035(.A1(n945), .A2(n935), .ZN(n1099));
  OAI22_X1  g1036(.A1(n939), .A2(n940), .B1(n794), .B2(n786), .ZN(n1100));
  INV_X1    g1037(.A(n934), .ZN(n1101));
  AOI21_X1  g1038(.A(n1101), .B1(n1093), .B2(n1091), .ZN(n1102));
  AND3_X1   g1039(.A1(n1101), .A2(n1093), .A3(n1091), .ZN(n1103));
  OAI221_X1 g1040(.A(n1100), .B1(n797), .B2(n796), .C1(n1103), .C2(n1102), .ZN(n1104));
  NAND3_X1  g1041(.A1(n1101), .A2(n1093), .A3(n1091), .ZN(n1105));
  OAI221_X1 g1042(.A(n1105), .B1(n933), .B2(n1094), .C1(n944), .C2(n936), .ZN(n1106));
  AOI21_X1  g1043(.A(n947), .B1(n1106), .B2(n1104), .ZN(n1107));
  NOR2_X1   g1044(.A1(n1107), .A2(n1099), .ZN(n1108));
  XNOR2_X1  g1045(.A(n1108), .B(n1098), .ZN(n1109));
  AND2_X1   g1046(.A1(426), .A2(103), .ZN(n1110));
  XNOR2_X1  g1047(.A(n1110), .B(n1109), .ZN(n1111));
  NOR2_X1   g1048(.A1(n958), .A2(n948), .ZN(n1112));
  OAI22_X1  g1049(.A1(n952), .A2(n953), .B1(n807), .B2(n799), .ZN(n1113));
  INV_X1    g1050(.A(n947), .ZN(n1114));
  AOI21_X1  g1051(.A(n1114), .B1(n1106), .B2(n1104), .ZN(n1115));
  AND3_X1   g1052(.A1(n1114), .A2(n1106), .A3(n1104), .ZN(n1116));
  OAI221_X1 g1053(.A(n1113), .B1(n810), .B2(n809), .C1(n1116), .C2(n1115), .ZN(n1117));
  NAND3_X1  g1054(.A1(n1114), .A2(n1106), .A3(n1104), .ZN(n1118));
  OAI221_X1 g1055(.A(n1118), .B1(n946), .B2(n1107), .C1(n957), .C2(n949), .ZN(n1119));
  AOI21_X1  g1056(.A(n960), .B1(n1119), .B2(n1117), .ZN(n1120));
  NOR2_X1   g1057(.A1(n1120), .A2(n1112), .ZN(n1121));
  XNOR2_X1  g1058(.A(n1121), .B(n1111), .ZN(n1122));
  AND2_X1   g1059(.A1(443), .A2(86), .ZN(n1123));
  XNOR2_X1  g1060(.A(n1123), .B(n1122), .ZN(n1124));
  NOR2_X1   g1061(.A1(n971), .A2(n961), .ZN(n1125));
  OAI22_X1  g1062(.A1(n965), .A2(n966), .B1(n820), .B2(n812), .ZN(n1126));
  INV_X1    g1063(.A(n960), .ZN(n1127));
  AOI21_X1  g1064(.A(n1127), .B1(n1119), .B2(n1117), .ZN(n1128));
  AND3_X1   g1065(.A1(n1127), .A2(n1119), .A3(n1117), .ZN(n1129));
  OAI221_X1 g1066(.A(n1126), .B1(n823), .B2(n822), .C1(n1129), .C2(n1128), .ZN(n1130));
  NAND3_X1  g1067(.A1(n1127), .A2(n1119), .A3(n1117), .ZN(n1131));
  OAI221_X1 g1068(.A(n1131), .B1(n959), .B2(n1120), .C1(n970), .C2(n962), .ZN(n1132));
  AOI21_X1  g1069(.A(n973), .B1(n1132), .B2(n1130), .ZN(n1133));
  NOR2_X1   g1070(.A1(n1133), .A2(n1125), .ZN(n1134));
  XNOR2_X1  g1071(.A(n1134), .B(n1124), .ZN(n1135));
  AND2_X1   g1072(.A1(460), .A2(69), .ZN(n1136));
  XNOR2_X1  g1073(.A(n1136), .B(n1135), .ZN(n1137));
  NOR2_X1   g1074(.A1(n984), .A2(n974), .ZN(n1138));
  OAI22_X1  g1075(.A1(n978), .A2(n979), .B1(n833), .B2(n825), .ZN(n1139));
  INV_X1    g1076(.A(n973), .ZN(n1140));
  AOI21_X1  g1077(.A(n1140), .B1(n1132), .B2(n1130), .ZN(n1141));
  AND3_X1   g1078(.A1(n1140), .A2(n1132), .A3(n1130), .ZN(n1142));
  OAI221_X1 g1079(.A(n1139), .B1(n836), .B2(n835), .C1(n1142), .C2(n1141), .ZN(n1143));
  NAND3_X1  g1080(.A1(n1140), .A2(n1132), .A3(n1130), .ZN(n1144));
  OAI221_X1 g1081(.A(n1144), .B1(n972), .B2(n1133), .C1(n983), .C2(n975), .ZN(n1145));
  AOI21_X1  g1082(.A(n986), .B1(n1145), .B2(n1143), .ZN(n1146));
  NOR2_X1   g1083(.A1(n1146), .A2(n1138), .ZN(n1147));
  XNOR2_X1  g1084(.A(n1147), .B(n1137), .ZN(n1148));
  AND2_X1   g1085(.A1(477), .A2(52), .ZN(n1149));
  XNOR2_X1  g1086(.A(n1149), .B(n1148), .ZN(n1150));
  NOR2_X1   g1087(.A1(n997), .A2(n987), .ZN(n1151));
  OAI22_X1  g1088(.A1(n991), .A2(n992), .B1(n846), .B2(n838), .ZN(n1152));
  INV_X1    g1089(.A(n986), .ZN(n1153));
  AOI21_X1  g1090(.A(n1153), .B1(n1145), .B2(n1143), .ZN(n1154));
  AND3_X1   g1091(.A1(n1153), .A2(n1145), .A3(n1143), .ZN(n1155));
  OAI221_X1 g1092(.A(n1152), .B1(n849), .B2(n848), .C1(n1155), .C2(n1154), .ZN(n1156));
  NAND3_X1  g1093(.A1(n1153), .A2(n1145), .A3(n1143), .ZN(n1157));
  OAI221_X1 g1094(.A(n1157), .B1(n985), .B2(n1146), .C1(n996), .C2(n988), .ZN(n1158));
  AOI21_X1  g1095(.A(n999), .B1(n1158), .B2(n1156), .ZN(n1159));
  NOR2_X1   g1096(.A1(n1159), .A2(n1151), .ZN(n1160));
  XNOR2_X1  g1097(.A(n1160), .B(n1150), .ZN(n1161));
  AND2_X1   g1098(.A1(494), .A2(35), .ZN(n1162));
  XNOR2_X1  g1099(.A(n1162), .B(n1161), .ZN(n1163));
  NOR2_X1   g1100(.A1(n1010), .A2(n1000), .ZN(n1164));
  OAI22_X1  g1101(.A1(n1004), .A2(n1005), .B1(n859), .B2(n851), .ZN(n1165));
  INV_X1    g1102(.A(n999), .ZN(n1166));
  AOI21_X1  g1103(.A(n1166), .B1(n1158), .B2(n1156), .ZN(n1167));
  AND3_X1   g1104(.A1(n1166), .A2(n1158), .A3(n1156), .ZN(n1168));
  OAI221_X1 g1105(.A(n1165), .B1(n862), .B2(n861), .C1(n1168), .C2(n1167), .ZN(n1169));
  NAND3_X1  g1106(.A1(n1166), .A2(n1158), .A3(n1156), .ZN(n1170));
  OAI221_X1 g1107(.A(n1170), .B1(n998), .B2(n1159), .C1(n1009), .C2(n1001), .ZN(n1171));
  AOI21_X1  g1108(.A(n1012), .B1(n1171), .B2(n1169), .ZN(n1172));
  NOR2_X1   g1109(.A1(n1172), .A2(n1164), .ZN(n1173));
  XNOR2_X1  g1110(.A(n1173), .B(n1163), .ZN(n1174));
  AND2_X1   g1111(.A1(511), .A2(18), .ZN(n1175));
  XNOR2_X1  g1112(.A(n1175), .B(n1174), .ZN(n1176));
  NOR2_X1   g1113(.A1(n1015), .A2(n1013), .ZN(n1177));
  AOI21_X1  g1114(.A(n1177), .B1(n1018), .B2(n1016), .ZN(n1178));
  XOR2_X1   g1115(.A(n1178), .B(n1176), .ZN(n1179));
  AND2_X1   g1116(.A1(528), .A2(\1 ), .ZN(n1180));
  INV_X1    g1117(.A(n1180), .ZN(n1181));
  XNOR2_X1  g1118(.A(n1181), .B(n1179), .ZN(6123));
  AND2_X1   g1119(.A1(290), .A2(256), .ZN(n1183));
  XOR2_X1   g1120(.A(n1183), .B(n1020), .ZN(n1184));
  NAND2_X1  g1121(.A1(307), .A2(239), .ZN(n1185));
  XNOR2_X1  g1122(.A(n1185), .B(n1184), .ZN(n1186));
  NOR2_X1   g1123(.A1(n1022), .A2(n870), .ZN(n1187));
  OAI21_X1  g1124(.A(n870), .B1(n1021), .B2(n1020), .ZN(n1188));
  OR3_X1    g1125(.A1(n1021), .A2(n1020), .A3(n870), .ZN(n1189));
  AOI21_X1  g1126(.A(n1024), .B1(n1189), .B2(n1188), .ZN(n1190));
  NOR2_X1   g1127(.A1(n1190), .A2(n1187), .ZN(n1191));
  XNOR2_X1  g1128(.A(n1191), .B(n1186), .ZN(n1192));
  AND2_X1   g1129(.A1(324), .A2(222), .ZN(n1193));
  XNOR2_X1  g1130(.A(n1193), .B(n1192), .ZN(n1194));
  NOR2_X1   g1131(.A1(n1030), .A2(n1025), .ZN(n1195));
  OR2_X1    g1132(.A1(n872), .A2(n733), .ZN(n1196));
  NAND2_X1  g1133(.A1(307), .A2(222), .ZN(n1197));
  AOI21_X1  g1134(.A(n1197), .B1(n1189), .B2(n1188), .ZN(n1198));
  AND3_X1   g1135(.A1(n1197), .A2(n1189), .A3(n1188), .ZN(n1199));
  OAI221_X1 g1136(.A(n1196), .B1(n874), .B2(n873), .C1(n1199), .C2(n1198), .ZN(n1200));
  NAND3_X1  g1137(.A1(n1197), .A2(n1189), .A3(n1188), .ZN(n1201));
  OAI221_X1 g1138(.A(n1201), .B1(n1023), .B2(n1190), .C1(n1029), .C2(n1026), .ZN(n1202));
  AOI21_X1  g1139(.A(n1032), .B1(n1202), .B2(n1200), .ZN(n1203));
  NOR2_X1   g1140(.A1(n1203), .A2(n1195), .ZN(n1204));
  XNOR2_X1  g1141(.A(n1204), .B(n1194), .ZN(n1205));
  AND2_X1   g1142(.A1(341), .A2(205), .ZN(n1206));
  XNOR2_X1  g1143(.A(n1206), .B(n1205), .ZN(n1207));
  NOR2_X1   g1144(.A1(n1043), .A2(n1033), .ZN(n1208));
  OAI22_X1  g1145(.A1(n1037), .A2(n1038), .B1(n879), .B2(n876), .ZN(n1209));
  INV_X1    g1146(.A(n1032), .ZN(n1210));
  AOI21_X1  g1147(.A(n1210), .B1(n1202), .B2(n1200), .ZN(n1211));
  AND3_X1   g1148(.A1(n1210), .A2(n1202), .A3(n1200), .ZN(n1212));
  OAI221_X1 g1149(.A(n1209), .B1(n882), .B2(n881), .C1(n1212), .C2(n1211), .ZN(n1213));
  NAND3_X1  g1150(.A1(n1210), .A2(n1202), .A3(n1200), .ZN(n1214));
  OAI221_X1 g1151(.A(n1214), .B1(n1031), .B2(n1203), .C1(n1042), .C2(n1034), .ZN(n1215));
  AOI21_X1  g1152(.A(n1045), .B1(n1215), .B2(n1213), .ZN(n1216));
  NOR2_X1   g1153(.A1(n1216), .A2(n1208), .ZN(n1217));
  XNOR2_X1  g1154(.A(n1217), .B(n1207), .ZN(n1218));
  AND2_X1   g1155(.A1(358), .A2(188), .ZN(n1219));
  XNOR2_X1  g1156(.A(n1219), .B(n1218), .ZN(n1220));
  NOR2_X1   g1157(.A1(n1056), .A2(n1046), .ZN(n1221));
  OAI22_X1  g1158(.A1(n1050), .A2(n1051), .B1(n892), .B2(n884), .ZN(n1222));
  INV_X1    g1159(.A(n1045), .ZN(n1223));
  AOI21_X1  g1160(.A(n1223), .B1(n1215), .B2(n1213), .ZN(n1224));
  AND3_X1   g1161(.A1(n1223), .A2(n1215), .A3(n1213), .ZN(n1225));
  OAI221_X1 g1162(.A(n1222), .B1(n895), .B2(n894), .C1(n1225), .C2(n1224), .ZN(n1226));
  NAND3_X1  g1163(.A1(n1223), .A2(n1215), .A3(n1213), .ZN(n1227));
  OAI221_X1 g1164(.A(n1227), .B1(n1044), .B2(n1216), .C1(n1055), .C2(n1047), .ZN(n1228));
  AOI21_X1  g1165(.A(n1058), .B1(n1228), .B2(n1226), .ZN(n1229));
  NOR2_X1   g1166(.A1(n1229), .A2(n1221), .ZN(n1230));
  XNOR2_X1  g1167(.A(n1230), .B(n1220), .ZN(n1231));
  AND2_X1   g1168(.A1(375), .A2(171), .ZN(n1232));
  XNOR2_X1  g1169(.A(n1232), .B(n1231), .ZN(n1233));
  NOR2_X1   g1170(.A1(n1069), .A2(n1059), .ZN(n1234));
  OAI22_X1  g1171(.A1(n1063), .A2(n1064), .B1(n905), .B2(n897), .ZN(n1235));
  INV_X1    g1172(.A(n1058), .ZN(n1236));
  AOI21_X1  g1173(.A(n1236), .B1(n1228), .B2(n1226), .ZN(n1237));
  AND3_X1   g1174(.A1(n1236), .A2(n1228), .A3(n1226), .ZN(n1238));
  OAI221_X1 g1175(.A(n1235), .B1(n908), .B2(n907), .C1(n1238), .C2(n1237), .ZN(n1239));
  NAND3_X1  g1176(.A1(n1236), .A2(n1228), .A3(n1226), .ZN(n1240));
  OAI221_X1 g1177(.A(n1240), .B1(n1057), .B2(n1229), .C1(n1068), .C2(n1060), .ZN(n1241));
  AOI21_X1  g1178(.A(n1071), .B1(n1241), .B2(n1239), .ZN(n1242));
  NOR2_X1   g1179(.A1(n1242), .A2(n1234), .ZN(n1243));
  XNOR2_X1  g1180(.A(n1243), .B(n1233), .ZN(n1244));
  AND2_X1   g1181(.A1(392), .A2(154), .ZN(n1245));
  XNOR2_X1  g1182(.A(n1245), .B(n1244), .ZN(n1246));
  NOR2_X1   g1183(.A1(n1082), .A2(n1072), .ZN(n1247));
  OAI22_X1  g1184(.A1(n1076), .A2(n1077), .B1(n918), .B2(n910), .ZN(n1248));
  INV_X1    g1185(.A(n1071), .ZN(n1249));
  AOI21_X1  g1186(.A(n1249), .B1(n1241), .B2(n1239), .ZN(n1250));
  AND3_X1   g1187(.A1(n1249), .A2(n1241), .A3(n1239), .ZN(n1251));
  OAI221_X1 g1188(.A(n1248), .B1(n921), .B2(n920), .C1(n1251), .C2(n1250), .ZN(n1252));
  NAND3_X1  g1189(.A1(n1249), .A2(n1241), .A3(n1239), .ZN(n1253));
  OAI221_X1 g1190(.A(n1253), .B1(n1070), .B2(n1242), .C1(n1081), .C2(n1073), .ZN(n1254));
  AOI21_X1  g1191(.A(n1084), .B1(n1254), .B2(n1252), .ZN(n1255));
  NOR2_X1   g1192(.A1(n1255), .A2(n1247), .ZN(n1256));
  XNOR2_X1  g1193(.A(n1256), .B(n1246), .ZN(n1257));
  AND2_X1   g1194(.A1(409), .A2(137), .ZN(n1258));
  XNOR2_X1  g1195(.A(n1258), .B(n1257), .ZN(n1259));
  NOR2_X1   g1196(.A1(n1095), .A2(n1085), .ZN(n1260));
  OAI22_X1  g1197(.A1(n1089), .A2(n1090), .B1(n931), .B2(n923), .ZN(n1261));
  INV_X1    g1198(.A(n1084), .ZN(n1262));
  AOI21_X1  g1199(.A(n1262), .B1(n1254), .B2(n1252), .ZN(n1263));
  AND3_X1   g1200(.A1(n1262), .A2(n1254), .A3(n1252), .ZN(n1264));
  OAI221_X1 g1201(.A(n1261), .B1(n934), .B2(n933), .C1(n1264), .C2(n1263), .ZN(n1265));
  NAND3_X1  g1202(.A1(n1262), .A2(n1254), .A3(n1252), .ZN(n1266));
  OAI221_X1 g1203(.A(n1266), .B1(n1083), .B2(n1255), .C1(n1094), .C2(n1086), .ZN(n1267));
  AOI21_X1  g1204(.A(n1097), .B1(n1267), .B2(n1265), .ZN(n1268));
  NOR2_X1   g1205(.A1(n1268), .A2(n1260), .ZN(n1269));
  XNOR2_X1  g1206(.A(n1269), .B(n1259), .ZN(n1270));
  AND2_X1   g1207(.A1(426), .A2(120), .ZN(n1271));
  XNOR2_X1  g1208(.A(n1271), .B(n1270), .ZN(n1272));
  NOR2_X1   g1209(.A1(n1108), .A2(n1098), .ZN(n1273));
  OAI22_X1  g1210(.A1(n1102), .A2(n1103), .B1(n944), .B2(n936), .ZN(n1274));
  INV_X1    g1211(.A(n1097), .ZN(n1275));
  AOI21_X1  g1212(.A(n1275), .B1(n1267), .B2(n1265), .ZN(n1276));
  AND3_X1   g1213(.A1(n1275), .A2(n1267), .A3(n1265), .ZN(n1277));
  OAI221_X1 g1214(.A(n1274), .B1(n947), .B2(n946), .C1(n1277), .C2(n1276), .ZN(n1278));
  NAND3_X1  g1215(.A1(n1275), .A2(n1267), .A3(n1265), .ZN(n1279));
  OAI221_X1 g1216(.A(n1279), .B1(n1096), .B2(n1268), .C1(n1107), .C2(n1099), .ZN(n1280));
  AOI21_X1  g1217(.A(n1110), .B1(n1280), .B2(n1278), .ZN(n1281));
  NOR2_X1   g1218(.A1(n1281), .A2(n1273), .ZN(n1282));
  XNOR2_X1  g1219(.A(n1282), .B(n1272), .ZN(n1283));
  AND2_X1   g1220(.A1(443), .A2(103), .ZN(n1284));
  XNOR2_X1  g1221(.A(n1284), .B(n1283), .ZN(n1285));
  NOR2_X1   g1222(.A1(n1121), .A2(n1111), .ZN(n1286));
  OAI22_X1  g1223(.A1(n1115), .A2(n1116), .B1(n957), .B2(n949), .ZN(n1287));
  INV_X1    g1224(.A(n1110), .ZN(n1288));
  AOI21_X1  g1225(.A(n1288), .B1(n1280), .B2(n1278), .ZN(n1289));
  AND3_X1   g1226(.A1(n1288), .A2(n1280), .A3(n1278), .ZN(n1290));
  OAI221_X1 g1227(.A(n1287), .B1(n960), .B2(n959), .C1(n1290), .C2(n1289), .ZN(n1291));
  NAND3_X1  g1228(.A1(n1288), .A2(n1280), .A3(n1278), .ZN(n1292));
  OAI221_X1 g1229(.A(n1292), .B1(n1109), .B2(n1281), .C1(n1120), .C2(n1112), .ZN(n1293));
  AOI21_X1  g1230(.A(n1123), .B1(n1293), .B2(n1291), .ZN(n1294));
  NOR2_X1   g1231(.A1(n1294), .A2(n1286), .ZN(n1295));
  XNOR2_X1  g1232(.A(n1295), .B(n1285), .ZN(n1296));
  AND2_X1   g1233(.A1(460), .A2(86), .ZN(n1297));
  XNOR2_X1  g1234(.A(n1297), .B(n1296), .ZN(n1298));
  NOR2_X1   g1235(.A1(n1134), .A2(n1124), .ZN(n1299));
  OAI22_X1  g1236(.A1(n1128), .A2(n1129), .B1(n970), .B2(n962), .ZN(n1300));
  INV_X1    g1237(.A(n1123), .ZN(n1301));
  AOI21_X1  g1238(.A(n1301), .B1(n1293), .B2(n1291), .ZN(n1302));
  AND3_X1   g1239(.A1(n1301), .A2(n1293), .A3(n1291), .ZN(n1303));
  OAI221_X1 g1240(.A(n1300), .B1(n973), .B2(n972), .C1(n1303), .C2(n1302), .ZN(n1304));
  NAND3_X1  g1241(.A1(n1301), .A2(n1293), .A3(n1291), .ZN(n1305));
  OAI221_X1 g1242(.A(n1305), .B1(n1122), .B2(n1294), .C1(n1133), .C2(n1125), .ZN(n1306));
  AOI21_X1  g1243(.A(n1136), .B1(n1306), .B2(n1304), .ZN(n1307));
  NOR2_X1   g1244(.A1(n1307), .A2(n1299), .ZN(n1308));
  XNOR2_X1  g1245(.A(n1308), .B(n1298), .ZN(n1309));
  AND2_X1   g1246(.A1(477), .A2(69), .ZN(n1310));
  XNOR2_X1  g1247(.A(n1310), .B(n1309), .ZN(n1311));
  NOR2_X1   g1248(.A1(n1147), .A2(n1137), .ZN(n1312));
  OAI22_X1  g1249(.A1(n1141), .A2(n1142), .B1(n983), .B2(n975), .ZN(n1313));
  INV_X1    g1250(.A(n1136), .ZN(n1314));
  AOI21_X1  g1251(.A(n1314), .B1(n1306), .B2(n1304), .ZN(n1315));
  AND3_X1   g1252(.A1(n1314), .A2(n1306), .A3(n1304), .ZN(n1316));
  OAI221_X1 g1253(.A(n1313), .B1(n986), .B2(n985), .C1(n1316), .C2(n1315), .ZN(n1317));
  NAND3_X1  g1254(.A1(n1314), .A2(n1306), .A3(n1304), .ZN(n1318));
  OAI221_X1 g1255(.A(n1318), .B1(n1135), .B2(n1307), .C1(n1146), .C2(n1138), .ZN(n1319));
  AOI21_X1  g1256(.A(n1149), .B1(n1319), .B2(n1317), .ZN(n1320));
  NOR2_X1   g1257(.A1(n1320), .A2(n1312), .ZN(n1321));
  XNOR2_X1  g1258(.A(n1321), .B(n1311), .ZN(n1322));
  AND2_X1   g1259(.A1(494), .A2(52), .ZN(n1323));
  XNOR2_X1  g1260(.A(n1323), .B(n1322), .ZN(n1324));
  NOR2_X1   g1261(.A1(n1160), .A2(n1150), .ZN(n1325));
  OAI22_X1  g1262(.A1(n1154), .A2(n1155), .B1(n996), .B2(n988), .ZN(n1326));
  INV_X1    g1263(.A(n1149), .ZN(n1327));
  AOI21_X1  g1264(.A(n1327), .B1(n1319), .B2(n1317), .ZN(n1328));
  AND3_X1   g1265(.A1(n1327), .A2(n1319), .A3(n1317), .ZN(n1329));
  OAI221_X1 g1266(.A(n1326), .B1(n999), .B2(n998), .C1(n1329), .C2(n1328), .ZN(n1330));
  NAND3_X1  g1267(.A1(n1327), .A2(n1319), .A3(n1317), .ZN(n1331));
  OAI221_X1 g1268(.A(n1331), .B1(n1148), .B2(n1320), .C1(n1159), .C2(n1151), .ZN(n1332));
  AOI21_X1  g1269(.A(n1162), .B1(n1332), .B2(n1330), .ZN(n1333));
  NOR2_X1   g1270(.A1(n1333), .A2(n1325), .ZN(n1334));
  XNOR2_X1  g1271(.A(n1334), .B(n1324), .ZN(n1335));
  AND2_X1   g1272(.A1(511), .A2(35), .ZN(n1336));
  XNOR2_X1  g1273(.A(n1336), .B(n1335), .ZN(n1337));
  NOR2_X1   g1274(.A1(n1173), .A2(n1163), .ZN(n1338));
  OAI22_X1  g1275(.A1(n1167), .A2(n1168), .B1(n1009), .B2(n1001), .ZN(n1339));
  INV_X1    g1276(.A(n1162), .ZN(n1340));
  AOI21_X1  g1277(.A(n1340), .B1(n1332), .B2(n1330), .ZN(n1341));
  AND3_X1   g1278(.A1(n1340), .A2(n1332), .A3(n1330), .ZN(n1342));
  OAI221_X1 g1279(.A(n1339), .B1(n1012), .B2(n1011), .C1(n1342), .C2(n1341), .ZN(n1343));
  NAND3_X1  g1280(.A1(n1340), .A2(n1332), .A3(n1330), .ZN(n1344));
  OAI221_X1 g1281(.A(n1344), .B1(n1161), .B2(n1333), .C1(n1172), .C2(n1164), .ZN(n1345));
  AOI21_X1  g1282(.A(n1175), .B1(n1345), .B2(n1343), .ZN(n1346));
  NOR2_X1   g1283(.A1(n1346), .A2(n1338), .ZN(n1347));
  XNOR2_X1  g1284(.A(n1347), .B(n1337), .ZN(n1348));
  AND2_X1   g1285(.A1(528), .A2(18), .ZN(n1349));
  XNOR2_X1  g1286(.A(n1349), .B(n1348), .ZN(n1350));
  NOR2_X1   g1287(.A1(n1178), .A2(n1176), .ZN(n1351));
  AOI21_X1  g1288(.A(n1351), .B1(n1181), .B2(n1179), .ZN(n1352));
  XOR2_X1   g1289(.A(n1352), .B(n1350), .ZN(6150));
  AND2_X1   g1290(.A1(307), .A2(256), .ZN(n1354));
  NOR2_X1   g1291(.A1(n1183), .A2(n1020), .ZN(n1355));
  AOI21_X1  g1292(.A(n1355), .B1(n1185), .B2(n1184), .ZN(n1356));
  XNOR2_X1  g1293(.A(n1356), .B(n1354), .ZN(n1357));
  AND2_X1   g1294(.A1(324), .A2(239), .ZN(n1358));
  XNOR2_X1  g1295(.A(n1358), .B(n1357), .ZN(n1359));
  NOR2_X1   g1296(.A1(n1191), .A2(n1186), .ZN(n1360));
  OR3_X1    g1297(.A1(n1186), .A2(n1190), .A3(n1187), .ZN(n1361));
  OAI21_X1  g1298(.A(n1186), .B1(n1190), .B2(n1187), .ZN(n1362));
  AOI21_X1  g1299(.A(n1193), .B1(n1362), .B2(n1361), .ZN(n1363));
  NOR2_X1   g1300(.A1(n1363), .A2(n1360), .ZN(n1364));
  XNOR2_X1  g1301(.A(n1364), .B(n1359), .ZN(n1365));
  AND2_X1   g1302(.A1(341), .A2(222), .ZN(n1366));
  XNOR2_X1  g1303(.A(n1366), .B(n1365), .ZN(n1367));
  NOR2_X1   g1304(.A1(n1204), .A2(n1194), .ZN(n1368));
  OAI22_X1  g1305(.A1(n1198), .A2(n1199), .B1(n1029), .B2(n1026), .ZN(n1369));
  INV_X1    g1306(.A(n1193), .ZN(n1370));
  AOI21_X1  g1307(.A(n1370), .B1(n1362), .B2(n1361), .ZN(n1371));
  AND3_X1   g1308(.A1(n1370), .A2(n1362), .A3(n1361), .ZN(n1372));
  OAI221_X1 g1309(.A(n1369), .B1(n1032), .B2(n1031), .C1(n1372), .C2(n1371), .ZN(n1373));
  NAND3_X1  g1310(.A1(n1370), .A2(n1362), .A3(n1361), .ZN(n1374));
  OAI221_X1 g1311(.A(n1374), .B1(n1192), .B2(n1363), .C1(n1203), .C2(n1195), .ZN(n1375));
  AOI21_X1  g1312(.A(n1206), .B1(n1375), .B2(n1373), .ZN(n1376));
  NOR2_X1   g1313(.A1(n1376), .A2(n1368), .ZN(n1377));
  XNOR2_X1  g1314(.A(n1377), .B(n1367), .ZN(n1378));
  AND2_X1   g1315(.A1(358), .A2(205), .ZN(n1379));
  XNOR2_X1  g1316(.A(n1379), .B(n1378), .ZN(n1380));
  NOR2_X1   g1317(.A1(n1217), .A2(n1207), .ZN(n1381));
  OAI22_X1  g1318(.A1(n1211), .A2(n1212), .B1(n1042), .B2(n1034), .ZN(n1382));
  INV_X1    g1319(.A(n1206), .ZN(n1383));
  AOI21_X1  g1320(.A(n1383), .B1(n1375), .B2(n1373), .ZN(n1384));
  AND3_X1   g1321(.A1(n1383), .A2(n1375), .A3(n1373), .ZN(n1385));
  OAI221_X1 g1322(.A(n1382), .B1(n1045), .B2(n1044), .C1(n1385), .C2(n1384), .ZN(n1386));
  NAND3_X1  g1323(.A1(n1383), .A2(n1375), .A3(n1373), .ZN(n1387));
  OAI221_X1 g1324(.A(n1387), .B1(n1205), .B2(n1376), .C1(n1216), .C2(n1208), .ZN(n1388));
  AOI21_X1  g1325(.A(n1219), .B1(n1388), .B2(n1386), .ZN(n1389));
  NOR2_X1   g1326(.A1(n1389), .A2(n1381), .ZN(n1390));
  XNOR2_X1  g1327(.A(n1390), .B(n1380), .ZN(n1391));
  AND2_X1   g1328(.A1(375), .A2(188), .ZN(n1392));
  XNOR2_X1  g1329(.A(n1392), .B(n1391), .ZN(n1393));
  NOR2_X1   g1330(.A1(n1230), .A2(n1220), .ZN(n1394));
  OAI22_X1  g1331(.A1(n1224), .A2(n1225), .B1(n1055), .B2(n1047), .ZN(n1395));
  INV_X1    g1332(.A(n1219), .ZN(n1396));
  AOI21_X1  g1333(.A(n1396), .B1(n1388), .B2(n1386), .ZN(n1397));
  AND3_X1   g1334(.A1(n1396), .A2(n1388), .A3(n1386), .ZN(n1398));
  OAI221_X1 g1335(.A(n1395), .B1(n1058), .B2(n1057), .C1(n1398), .C2(n1397), .ZN(n1399));
  NAND3_X1  g1336(.A1(n1396), .A2(n1388), .A3(n1386), .ZN(n1400));
  OAI221_X1 g1337(.A(n1400), .B1(n1218), .B2(n1389), .C1(n1229), .C2(n1221), .ZN(n1401));
  AOI21_X1  g1338(.A(n1232), .B1(n1401), .B2(n1399), .ZN(n1402));
  NOR2_X1   g1339(.A1(n1402), .A2(n1394), .ZN(n1403));
  XNOR2_X1  g1340(.A(n1403), .B(n1393), .ZN(n1404));
  AND2_X1   g1341(.A1(392), .A2(171), .ZN(n1405));
  XNOR2_X1  g1342(.A(n1405), .B(n1404), .ZN(n1406));
  NOR2_X1   g1343(.A1(n1243), .A2(n1233), .ZN(n1407));
  OAI22_X1  g1344(.A1(n1237), .A2(n1238), .B1(n1068), .B2(n1060), .ZN(n1408));
  INV_X1    g1345(.A(n1232), .ZN(n1409));
  AOI21_X1  g1346(.A(n1409), .B1(n1401), .B2(n1399), .ZN(n1410));
  AND3_X1   g1347(.A1(n1409), .A2(n1401), .A3(n1399), .ZN(n1411));
  OAI221_X1 g1348(.A(n1408), .B1(n1071), .B2(n1070), .C1(n1411), .C2(n1410), .ZN(n1412));
  NAND3_X1  g1349(.A1(n1409), .A2(n1401), .A3(n1399), .ZN(n1413));
  OAI221_X1 g1350(.A(n1413), .B1(n1231), .B2(n1402), .C1(n1242), .C2(n1234), .ZN(n1414));
  AOI21_X1  g1351(.A(n1245), .B1(n1414), .B2(n1412), .ZN(n1415));
  NOR2_X1   g1352(.A1(n1415), .A2(n1407), .ZN(n1416));
  XNOR2_X1  g1353(.A(n1416), .B(n1406), .ZN(n1417));
  AND2_X1   g1354(.A1(409), .A2(154), .ZN(n1418));
  XNOR2_X1  g1355(.A(n1418), .B(n1417), .ZN(n1419));
  NOR2_X1   g1356(.A1(n1256), .A2(n1246), .ZN(n1420));
  OAI22_X1  g1357(.A1(n1250), .A2(n1251), .B1(n1081), .B2(n1073), .ZN(n1421));
  INV_X1    g1358(.A(n1245), .ZN(n1422));
  AOI21_X1  g1359(.A(n1422), .B1(n1414), .B2(n1412), .ZN(n1423));
  AND3_X1   g1360(.A1(n1422), .A2(n1414), .A3(n1412), .ZN(n1424));
  OAI221_X1 g1361(.A(n1421), .B1(n1084), .B2(n1083), .C1(n1424), .C2(n1423), .ZN(n1425));
  NAND3_X1  g1362(.A1(n1422), .A2(n1414), .A3(n1412), .ZN(n1426));
  OAI221_X1 g1363(.A(n1426), .B1(n1244), .B2(n1415), .C1(n1255), .C2(n1247), .ZN(n1427));
  AOI21_X1  g1364(.A(n1258), .B1(n1427), .B2(n1425), .ZN(n1428));
  NOR2_X1   g1365(.A1(n1428), .A2(n1420), .ZN(n1429));
  XNOR2_X1  g1366(.A(n1429), .B(n1419), .ZN(n1430));
  AND2_X1   g1367(.A1(426), .A2(137), .ZN(n1431));
  XNOR2_X1  g1368(.A(n1431), .B(n1430), .ZN(n1432));
  NOR2_X1   g1369(.A1(n1269), .A2(n1259), .ZN(n1433));
  OAI22_X1  g1370(.A1(n1263), .A2(n1264), .B1(n1094), .B2(n1086), .ZN(n1434));
  INV_X1    g1371(.A(n1258), .ZN(n1435));
  AOI21_X1  g1372(.A(n1435), .B1(n1427), .B2(n1425), .ZN(n1436));
  AND3_X1   g1373(.A1(n1435), .A2(n1427), .A3(n1425), .ZN(n1437));
  OAI221_X1 g1374(.A(n1434), .B1(n1097), .B2(n1096), .C1(n1437), .C2(n1436), .ZN(n1438));
  NAND3_X1  g1375(.A1(n1435), .A2(n1427), .A3(n1425), .ZN(n1439));
  OAI221_X1 g1376(.A(n1439), .B1(n1257), .B2(n1428), .C1(n1268), .C2(n1260), .ZN(n1440));
  AOI21_X1  g1377(.A(n1271), .B1(n1440), .B2(n1438), .ZN(n1441));
  NOR2_X1   g1378(.A1(n1441), .A2(n1433), .ZN(n1442));
  XNOR2_X1  g1379(.A(n1442), .B(n1432), .ZN(n1443));
  AND2_X1   g1380(.A1(443), .A2(120), .ZN(n1444));
  XNOR2_X1  g1381(.A(n1444), .B(n1443), .ZN(n1445));
  NOR2_X1   g1382(.A1(n1282), .A2(n1272), .ZN(n1446));
  OAI22_X1  g1383(.A1(n1276), .A2(n1277), .B1(n1107), .B2(n1099), .ZN(n1447));
  INV_X1    g1384(.A(n1271), .ZN(n1448));
  AOI21_X1  g1385(.A(n1448), .B1(n1440), .B2(n1438), .ZN(n1449));
  AND3_X1   g1386(.A1(n1448), .A2(n1440), .A3(n1438), .ZN(n1450));
  OAI221_X1 g1387(.A(n1447), .B1(n1110), .B2(n1109), .C1(n1450), .C2(n1449), .ZN(n1451));
  NAND3_X1  g1388(.A1(n1448), .A2(n1440), .A3(n1438), .ZN(n1452));
  OAI221_X1 g1389(.A(n1452), .B1(n1270), .B2(n1441), .C1(n1281), .C2(n1273), .ZN(n1453));
  AOI21_X1  g1390(.A(n1284), .B1(n1453), .B2(n1451), .ZN(n1454));
  NOR2_X1   g1391(.A1(n1454), .A2(n1446), .ZN(n1455));
  XNOR2_X1  g1392(.A(n1455), .B(n1445), .ZN(n1456));
  AND2_X1   g1393(.A1(460), .A2(103), .ZN(n1457));
  XNOR2_X1  g1394(.A(n1457), .B(n1456), .ZN(n1458));
  NOR2_X1   g1395(.A1(n1295), .A2(n1285), .ZN(n1459));
  OAI22_X1  g1396(.A1(n1289), .A2(n1290), .B1(n1120), .B2(n1112), .ZN(n1460));
  INV_X1    g1397(.A(n1284), .ZN(n1461));
  AOI21_X1  g1398(.A(n1461), .B1(n1453), .B2(n1451), .ZN(n1462));
  AND3_X1   g1399(.A1(n1461), .A2(n1453), .A3(n1451), .ZN(n1463));
  OAI221_X1 g1400(.A(n1460), .B1(n1123), .B2(n1122), .C1(n1463), .C2(n1462), .ZN(n1464));
  NAND3_X1  g1401(.A1(n1461), .A2(n1453), .A3(n1451), .ZN(n1465));
  OAI221_X1 g1402(.A(n1465), .B1(n1283), .B2(n1454), .C1(n1294), .C2(n1286), .ZN(n1466));
  AOI21_X1  g1403(.A(n1297), .B1(n1466), .B2(n1464), .ZN(n1467));
  NOR2_X1   g1404(.A1(n1467), .A2(n1459), .ZN(n1468));
  XNOR2_X1  g1405(.A(n1468), .B(n1458), .ZN(n1469));
  AND2_X1   g1406(.A1(477), .A2(86), .ZN(n1470));
  XNOR2_X1  g1407(.A(n1470), .B(n1469), .ZN(n1471));
  NOR2_X1   g1408(.A1(n1308), .A2(n1298), .ZN(n1472));
  OAI22_X1  g1409(.A1(n1302), .A2(n1303), .B1(n1133), .B2(n1125), .ZN(n1473));
  INV_X1    g1410(.A(n1297), .ZN(n1474));
  AOI21_X1  g1411(.A(n1474), .B1(n1466), .B2(n1464), .ZN(n1475));
  AND3_X1   g1412(.A1(n1474), .A2(n1466), .A3(n1464), .ZN(n1476));
  OAI221_X1 g1413(.A(n1473), .B1(n1136), .B2(n1135), .C1(n1476), .C2(n1475), .ZN(n1477));
  NAND3_X1  g1414(.A1(n1474), .A2(n1466), .A3(n1464), .ZN(n1478));
  OAI221_X1 g1415(.A(n1478), .B1(n1296), .B2(n1467), .C1(n1307), .C2(n1299), .ZN(n1479));
  AOI21_X1  g1416(.A(n1310), .B1(n1479), .B2(n1477), .ZN(n1480));
  NOR2_X1   g1417(.A1(n1480), .A2(n1472), .ZN(n1481));
  XNOR2_X1  g1418(.A(n1481), .B(n1471), .ZN(n1482));
  AND2_X1   g1419(.A1(494), .A2(69), .ZN(n1483));
  XNOR2_X1  g1420(.A(n1483), .B(n1482), .ZN(n1484));
  NOR2_X1   g1421(.A1(n1321), .A2(n1311), .ZN(n1485));
  OAI22_X1  g1422(.A1(n1315), .A2(n1316), .B1(n1146), .B2(n1138), .ZN(n1486));
  INV_X1    g1423(.A(n1310), .ZN(n1487));
  AOI21_X1  g1424(.A(n1487), .B1(n1479), .B2(n1477), .ZN(n1488));
  AND3_X1   g1425(.A1(n1487), .A2(n1479), .A3(n1477), .ZN(n1489));
  OAI221_X1 g1426(.A(n1486), .B1(n1149), .B2(n1148), .C1(n1489), .C2(n1488), .ZN(n1490));
  NAND3_X1  g1427(.A1(n1487), .A2(n1479), .A3(n1477), .ZN(n1491));
  OAI221_X1 g1428(.A(n1491), .B1(n1309), .B2(n1480), .C1(n1320), .C2(n1312), .ZN(n1492));
  AOI21_X1  g1429(.A(n1323), .B1(n1492), .B2(n1490), .ZN(n1493));
  NOR2_X1   g1430(.A1(n1493), .A2(n1485), .ZN(n1494));
  XNOR2_X1  g1431(.A(n1494), .B(n1484), .ZN(n1495));
  AND2_X1   g1432(.A1(511), .A2(52), .ZN(n1496));
  XNOR2_X1  g1433(.A(n1496), .B(n1495), .ZN(n1497));
  NOR2_X1   g1434(.A1(n1334), .A2(n1324), .ZN(n1498));
  OAI22_X1  g1435(.A1(n1328), .A2(n1329), .B1(n1159), .B2(n1151), .ZN(n1499));
  INV_X1    g1436(.A(n1323), .ZN(n1500));
  AOI21_X1  g1437(.A(n1500), .B1(n1492), .B2(n1490), .ZN(n1501));
  AND3_X1   g1438(.A1(n1500), .A2(n1492), .A3(n1490), .ZN(n1502));
  OAI221_X1 g1439(.A(n1499), .B1(n1162), .B2(n1161), .C1(n1502), .C2(n1501), .ZN(n1503));
  NAND3_X1  g1440(.A1(n1500), .A2(n1492), .A3(n1490), .ZN(n1504));
  OAI221_X1 g1441(.A(n1504), .B1(n1322), .B2(n1493), .C1(n1333), .C2(n1325), .ZN(n1505));
  AOI21_X1  g1442(.A(n1336), .B1(n1505), .B2(n1503), .ZN(n1506));
  NOR2_X1   g1443(.A1(n1506), .A2(n1498), .ZN(n1507));
  XNOR2_X1  g1444(.A(n1507), .B(n1497), .ZN(n1508));
  NAND2_X1  g1445(.A1(528), .A2(35), .ZN(n1509));
  XOR2_X1   g1446(.A(n1509), .B(n1508), .ZN(n1510));
  NOR2_X1   g1447(.A1(n1347), .A2(n1337), .ZN(n1511));
  OAI22_X1  g1448(.A1(n1341), .A2(n1342), .B1(n1172), .B2(n1164), .ZN(n1512));
  INV_X1    g1449(.A(n1336), .ZN(n1513));
  AOI21_X1  g1450(.A(n1513), .B1(n1505), .B2(n1503), .ZN(n1514));
  AND3_X1   g1451(.A1(n1513), .A2(n1505), .A3(n1503), .ZN(n1515));
  OAI221_X1 g1452(.A(n1512), .B1(n1175), .B2(n1174), .C1(n1515), .C2(n1514), .ZN(n1516));
  NAND3_X1  g1453(.A1(n1513), .A2(n1505), .A3(n1503), .ZN(n1517));
  OAI221_X1 g1454(.A(n1517), .B1(n1335), .B2(n1506), .C1(n1346), .C2(n1338), .ZN(n1518));
  AOI21_X1  g1455(.A(n1349), .B1(n1518), .B2(n1516), .ZN(n1519));
  NOR2_X1   g1456(.A1(n1519), .A2(n1511), .ZN(n1520));
  XNOR2_X1  g1457(.A(n1520), .B(n1510), .ZN(n1521));
  AND2_X1   g1458(.A1(n1352), .A2(n1350), .ZN(n1522));
  XNOR2_X1  g1459(.A(n1522), .B(n1521), .ZN(6160));
  AND2_X1   g1460(.A1(324), .A2(256), .ZN(n1524));
  NOR2_X1   g1461(.A1(n1356), .A2(n1354), .ZN(n1525));
  NOR2_X1   g1462(.A1(n1358), .A2(n1357), .ZN(n1526));
  NOR2_X1   g1463(.A1(n1526), .A2(n1525), .ZN(n1527));
  XNOR2_X1  g1464(.A(n1527), .B(n1524), .ZN(n1528));
  AND2_X1   g1465(.A1(341), .A2(239), .ZN(n1529));
  XNOR2_X1  g1466(.A(n1529), .B(n1528), .ZN(n1530));
  NOR2_X1   g1467(.A1(n1364), .A2(n1359), .ZN(n1531));
  OR3_X1    g1468(.A1(n1359), .A2(n1363), .A3(n1360), .ZN(n1532));
  OAI21_X1  g1469(.A(n1359), .B1(n1363), .B2(n1360), .ZN(n1533));
  AOI21_X1  g1470(.A(n1366), .B1(n1533), .B2(n1532), .ZN(n1534));
  NOR2_X1   g1471(.A1(n1534), .A2(n1531), .ZN(n1535));
  XNOR2_X1  g1472(.A(n1535), .B(n1530), .ZN(n1536));
  AND2_X1   g1473(.A1(358), .A2(222), .ZN(n1537));
  XNOR2_X1  g1474(.A(n1537), .B(n1536), .ZN(n1538));
  NOR2_X1   g1475(.A1(n1377), .A2(n1367), .ZN(n1539));
  OAI22_X1  g1476(.A1(n1371), .A2(n1372), .B1(n1203), .B2(n1195), .ZN(n1540));
  INV_X1    g1477(.A(n1366), .ZN(n1541));
  AOI21_X1  g1478(.A(n1541), .B1(n1533), .B2(n1532), .ZN(n1542));
  AND3_X1   g1479(.A1(n1541), .A2(n1533), .A3(n1532), .ZN(n1543));
  OAI221_X1 g1480(.A(n1540), .B1(n1206), .B2(n1205), .C1(n1543), .C2(n1542), .ZN(n1544));
  NAND3_X1  g1481(.A1(n1541), .A2(n1533), .A3(n1532), .ZN(n1545));
  OAI221_X1 g1482(.A(n1545), .B1(n1365), .B2(n1534), .C1(n1376), .C2(n1368), .ZN(n1546));
  AOI21_X1  g1483(.A(n1379), .B1(n1546), .B2(n1544), .ZN(n1547));
  NOR2_X1   g1484(.A1(n1547), .A2(n1539), .ZN(n1548));
  XNOR2_X1  g1485(.A(n1548), .B(n1538), .ZN(n1549));
  AND2_X1   g1486(.A1(375), .A2(205), .ZN(n1550));
  XNOR2_X1  g1487(.A(n1550), .B(n1549), .ZN(n1551));
  NOR2_X1   g1488(.A1(n1390), .A2(n1380), .ZN(n1552));
  OAI22_X1  g1489(.A1(n1384), .A2(n1385), .B1(n1216), .B2(n1208), .ZN(n1553));
  INV_X1    g1490(.A(n1379), .ZN(n1554));
  AOI21_X1  g1491(.A(n1554), .B1(n1546), .B2(n1544), .ZN(n1555));
  AND3_X1   g1492(.A1(n1554), .A2(n1546), .A3(n1544), .ZN(n1556));
  OAI221_X1 g1493(.A(n1553), .B1(n1219), .B2(n1218), .C1(n1556), .C2(n1555), .ZN(n1557));
  NAND3_X1  g1494(.A1(n1554), .A2(n1546), .A3(n1544), .ZN(n1558));
  OAI221_X1 g1495(.A(n1558), .B1(n1378), .B2(n1547), .C1(n1389), .C2(n1381), .ZN(n1559));
  AOI21_X1  g1496(.A(n1392), .B1(n1559), .B2(n1557), .ZN(n1560));
  NOR2_X1   g1497(.A1(n1560), .A2(n1552), .ZN(n1561));
  XNOR2_X1  g1498(.A(n1561), .B(n1551), .ZN(n1562));
  AND2_X1   g1499(.A1(392), .A2(188), .ZN(n1563));
  XNOR2_X1  g1500(.A(n1563), .B(n1562), .ZN(n1564));
  NOR2_X1   g1501(.A1(n1403), .A2(n1393), .ZN(n1565));
  OAI22_X1  g1502(.A1(n1397), .A2(n1398), .B1(n1229), .B2(n1221), .ZN(n1566));
  INV_X1    g1503(.A(n1392), .ZN(n1567));
  AOI21_X1  g1504(.A(n1567), .B1(n1559), .B2(n1557), .ZN(n1568));
  AND3_X1   g1505(.A1(n1567), .A2(n1559), .A3(n1557), .ZN(n1569));
  OAI221_X1 g1506(.A(n1566), .B1(n1232), .B2(n1231), .C1(n1569), .C2(n1568), .ZN(n1570));
  NAND3_X1  g1507(.A1(n1567), .A2(n1559), .A3(n1557), .ZN(n1571));
  OAI221_X1 g1508(.A(n1571), .B1(n1391), .B2(n1560), .C1(n1402), .C2(n1394), .ZN(n1572));
  AOI21_X1  g1509(.A(n1405), .B1(n1572), .B2(n1570), .ZN(n1573));
  NOR2_X1   g1510(.A1(n1573), .A2(n1565), .ZN(n1574));
  XNOR2_X1  g1511(.A(n1574), .B(n1564), .ZN(n1575));
  AND2_X1   g1512(.A1(409), .A2(171), .ZN(n1576));
  XNOR2_X1  g1513(.A(n1576), .B(n1575), .ZN(n1577));
  NOR2_X1   g1514(.A1(n1416), .A2(n1406), .ZN(n1578));
  OAI22_X1  g1515(.A1(n1410), .A2(n1411), .B1(n1242), .B2(n1234), .ZN(n1579));
  INV_X1    g1516(.A(n1405), .ZN(n1580));
  AOI21_X1  g1517(.A(n1580), .B1(n1572), .B2(n1570), .ZN(n1581));
  AND3_X1   g1518(.A1(n1580), .A2(n1572), .A3(n1570), .ZN(n1582));
  OAI221_X1 g1519(.A(n1579), .B1(n1245), .B2(n1244), .C1(n1582), .C2(n1581), .ZN(n1583));
  NAND3_X1  g1520(.A1(n1580), .A2(n1572), .A3(n1570), .ZN(n1584));
  OAI221_X1 g1521(.A(n1584), .B1(n1404), .B2(n1573), .C1(n1415), .C2(n1407), .ZN(n1585));
  AOI21_X1  g1522(.A(n1418), .B1(n1585), .B2(n1583), .ZN(n1586));
  NOR2_X1   g1523(.A1(n1586), .A2(n1578), .ZN(n1587));
  XNOR2_X1  g1524(.A(n1587), .B(n1577), .ZN(n1588));
  AND2_X1   g1525(.A1(426), .A2(154), .ZN(n1589));
  XNOR2_X1  g1526(.A(n1589), .B(n1588), .ZN(n1590));
  NOR2_X1   g1527(.A1(n1429), .A2(n1419), .ZN(n1591));
  OAI22_X1  g1528(.A1(n1423), .A2(n1424), .B1(n1255), .B2(n1247), .ZN(n1592));
  INV_X1    g1529(.A(n1418), .ZN(n1593));
  AOI21_X1  g1530(.A(n1593), .B1(n1585), .B2(n1583), .ZN(n1594));
  AND3_X1   g1531(.A1(n1593), .A2(n1585), .A3(n1583), .ZN(n1595));
  OAI221_X1 g1532(.A(n1592), .B1(n1258), .B2(n1257), .C1(n1595), .C2(n1594), .ZN(n1596));
  NAND3_X1  g1533(.A1(n1593), .A2(n1585), .A3(n1583), .ZN(n1597));
  OAI221_X1 g1534(.A(n1597), .B1(n1417), .B2(n1586), .C1(n1428), .C2(n1420), .ZN(n1598));
  AOI21_X1  g1535(.A(n1431), .B1(n1598), .B2(n1596), .ZN(n1599));
  NOR2_X1   g1536(.A1(n1599), .A2(n1591), .ZN(n1600));
  XNOR2_X1  g1537(.A(n1600), .B(n1590), .ZN(n1601));
  AND2_X1   g1538(.A1(443), .A2(137), .ZN(n1602));
  XNOR2_X1  g1539(.A(n1602), .B(n1601), .ZN(n1603));
  NOR2_X1   g1540(.A1(n1442), .A2(n1432), .ZN(n1604));
  OAI22_X1  g1541(.A1(n1436), .A2(n1437), .B1(n1268), .B2(n1260), .ZN(n1605));
  INV_X1    g1542(.A(n1431), .ZN(n1606));
  AOI21_X1  g1543(.A(n1606), .B1(n1598), .B2(n1596), .ZN(n1607));
  AND3_X1   g1544(.A1(n1606), .A2(n1598), .A3(n1596), .ZN(n1608));
  OAI221_X1 g1545(.A(n1605), .B1(n1271), .B2(n1270), .C1(n1608), .C2(n1607), .ZN(n1609));
  NAND3_X1  g1546(.A1(n1606), .A2(n1598), .A3(n1596), .ZN(n1610));
  OAI221_X1 g1547(.A(n1610), .B1(n1430), .B2(n1599), .C1(n1441), .C2(n1433), .ZN(n1611));
  AOI21_X1  g1548(.A(n1444), .B1(n1611), .B2(n1609), .ZN(n1612));
  NOR2_X1   g1549(.A1(n1612), .A2(n1604), .ZN(n1613));
  XNOR2_X1  g1550(.A(n1613), .B(n1603), .ZN(n1614));
  AND2_X1   g1551(.A1(460), .A2(120), .ZN(n1615));
  XNOR2_X1  g1552(.A(n1615), .B(n1614), .ZN(n1616));
  NOR2_X1   g1553(.A1(n1455), .A2(n1445), .ZN(n1617));
  OAI22_X1  g1554(.A1(n1449), .A2(n1450), .B1(n1281), .B2(n1273), .ZN(n1618));
  INV_X1    g1555(.A(n1444), .ZN(n1619));
  AOI21_X1  g1556(.A(n1619), .B1(n1611), .B2(n1609), .ZN(n1620));
  AND3_X1   g1557(.A1(n1619), .A2(n1611), .A3(n1609), .ZN(n1621));
  OAI221_X1 g1558(.A(n1618), .B1(n1284), .B2(n1283), .C1(n1621), .C2(n1620), .ZN(n1622));
  NAND3_X1  g1559(.A1(n1619), .A2(n1611), .A3(n1609), .ZN(n1623));
  OAI221_X1 g1560(.A(n1623), .B1(n1443), .B2(n1612), .C1(n1454), .C2(n1446), .ZN(n1624));
  AOI21_X1  g1561(.A(n1457), .B1(n1624), .B2(n1622), .ZN(n1625));
  NOR2_X1   g1562(.A1(n1625), .A2(n1617), .ZN(n1626));
  XNOR2_X1  g1563(.A(n1626), .B(n1616), .ZN(n1627));
  AND2_X1   g1564(.A1(477), .A2(103), .ZN(n1628));
  XNOR2_X1  g1565(.A(n1628), .B(n1627), .ZN(n1629));
  NOR2_X1   g1566(.A1(n1468), .A2(n1458), .ZN(n1630));
  OAI22_X1  g1567(.A1(n1462), .A2(n1463), .B1(n1294), .B2(n1286), .ZN(n1631));
  INV_X1    g1568(.A(n1457), .ZN(n1632));
  AOI21_X1  g1569(.A(n1632), .B1(n1624), .B2(n1622), .ZN(n1633));
  AND3_X1   g1570(.A1(n1632), .A2(n1624), .A3(n1622), .ZN(n1634));
  OAI221_X1 g1571(.A(n1631), .B1(n1297), .B2(n1296), .C1(n1634), .C2(n1633), .ZN(n1635));
  NAND3_X1  g1572(.A1(n1632), .A2(n1624), .A3(n1622), .ZN(n1636));
  OAI221_X1 g1573(.A(n1636), .B1(n1456), .B2(n1625), .C1(n1467), .C2(n1459), .ZN(n1637));
  AOI21_X1  g1574(.A(n1470), .B1(n1637), .B2(n1635), .ZN(n1638));
  NOR2_X1   g1575(.A1(n1638), .A2(n1630), .ZN(n1639));
  XNOR2_X1  g1576(.A(n1639), .B(n1629), .ZN(n1640));
  AND2_X1   g1577(.A1(494), .A2(86), .ZN(n1641));
  XNOR2_X1  g1578(.A(n1641), .B(n1640), .ZN(n1642));
  NOR2_X1   g1579(.A1(n1481), .A2(n1471), .ZN(n1643));
  OAI22_X1  g1580(.A1(n1475), .A2(n1476), .B1(n1307), .B2(n1299), .ZN(n1644));
  INV_X1    g1581(.A(n1470), .ZN(n1645));
  AOI21_X1  g1582(.A(n1645), .B1(n1637), .B2(n1635), .ZN(n1646));
  AND3_X1   g1583(.A1(n1645), .A2(n1637), .A3(n1635), .ZN(n1647));
  OAI221_X1 g1584(.A(n1644), .B1(n1310), .B2(n1309), .C1(n1647), .C2(n1646), .ZN(n1648));
  NAND3_X1  g1585(.A1(n1645), .A2(n1637), .A3(n1635), .ZN(n1649));
  OAI221_X1 g1586(.A(n1649), .B1(n1469), .B2(n1638), .C1(n1480), .C2(n1472), .ZN(n1650));
  AOI21_X1  g1587(.A(n1483), .B1(n1650), .B2(n1648), .ZN(n1651));
  NOR2_X1   g1588(.A1(n1651), .A2(n1643), .ZN(n1652));
  XNOR2_X1  g1589(.A(n1652), .B(n1642), .ZN(n1653));
  AND2_X1   g1590(.A1(511), .A2(69), .ZN(n1654));
  XNOR2_X1  g1591(.A(n1654), .B(n1653), .ZN(n1655));
  NOR2_X1   g1592(.A1(n1494), .A2(n1484), .ZN(n1656));
  OAI22_X1  g1593(.A1(n1488), .A2(n1489), .B1(n1320), .B2(n1312), .ZN(n1657));
  INV_X1    g1594(.A(n1483), .ZN(n1658));
  AOI21_X1  g1595(.A(n1658), .B1(n1650), .B2(n1648), .ZN(n1659));
  AND3_X1   g1596(.A1(n1658), .A2(n1650), .A3(n1648), .ZN(n1660));
  OAI221_X1 g1597(.A(n1657), .B1(n1323), .B2(n1322), .C1(n1660), .C2(n1659), .ZN(n1661));
  NAND3_X1  g1598(.A1(n1658), .A2(n1650), .A3(n1648), .ZN(n1662));
  OAI221_X1 g1599(.A(n1662), .B1(n1482), .B2(n1651), .C1(n1493), .C2(n1485), .ZN(n1663));
  AOI21_X1  g1600(.A(n1496), .B1(n1663), .B2(n1661), .ZN(n1664));
  NOR2_X1   g1601(.A1(n1664), .A2(n1656), .ZN(n1665));
  XOR2_X1   g1602(.A(n1665), .B(n1655), .ZN(n1666));
  NAND2_X1  g1603(.A1(528), .A2(52), .ZN(n1667));
  XNOR2_X1  g1604(.A(n1667), .B(n1666), .ZN(n1668));
  NOR2_X1   g1605(.A1(n1507), .A2(n1497), .ZN(n1669));
  OAI22_X1  g1606(.A1(n1501), .A2(n1502), .B1(n1333), .B2(n1325), .ZN(n1670));
  INV_X1    g1607(.A(n1496), .ZN(n1671));
  AOI21_X1  g1608(.A(n1671), .B1(n1663), .B2(n1661), .ZN(n1672));
  AND3_X1   g1609(.A1(n1671), .A2(n1663), .A3(n1661), .ZN(n1673));
  OAI221_X1 g1610(.A(n1670), .B1(n1336), .B2(n1335), .C1(n1673), .C2(n1672), .ZN(n1674));
  NAND3_X1  g1611(.A1(n1671), .A2(n1663), .A3(n1661), .ZN(n1675));
  OAI221_X1 g1612(.A(n1675), .B1(n1495), .B2(n1664), .C1(n1506), .C2(n1498), .ZN(n1676));
  AOI22_X1  g1613(.A1(n1674), .A2(n1676), .B1(528), .B2(35), .ZN(n1677));
  NOR2_X1   g1614(.A1(n1677), .A2(n1669), .ZN(n1678));
  XOR2_X1   g1615(.A(n1678), .B(n1668), .ZN(n1679));
  NOR2_X1   g1616(.A1(n1520), .A2(n1510), .ZN(n1680));
  OAI22_X1  g1617(.A1(n1514), .A2(n1515), .B1(n1346), .B2(n1338), .ZN(n1681));
  AOI21_X1  g1618(.A(n1509), .B1(n1676), .B2(n1674), .ZN(n1682));
  AND3_X1   g1619(.A1(n1509), .A2(n1676), .A3(n1674), .ZN(n1683));
  OAI221_X1 g1620(.A(n1681), .B1(n1349), .B2(n1348), .C1(n1683), .C2(n1682), .ZN(n1684));
  NAND3_X1  g1621(.A1(n1509), .A2(n1676), .A3(n1674), .ZN(n1685));
  OAI221_X1 g1622(.A(n1685), .B1(n1508), .B2(n1677), .C1(n1519), .C2(n1511), .ZN(n1686));
  AOI22_X1  g1623(.A1(n1684), .A2(n1686), .B1(n1352), .B2(n1350), .ZN(n1687));
  OR2_X1    g1624(.A1(n1687), .A2(n1680), .ZN(n1688));
  XNOR2_X1  g1625(.A(n1688), .B(n1679), .ZN(6170));
  AND2_X1   g1626(.A1(341), .A2(256), .ZN(n1690));
  NOR2_X1   g1627(.A1(n1527), .A2(n1524), .ZN(n1691));
  NOR2_X1   g1628(.A1(n1529), .A2(n1528), .ZN(n1692));
  NOR2_X1   g1629(.A1(n1692), .A2(n1691), .ZN(n1693));
  XNOR2_X1  g1630(.A(n1693), .B(n1690), .ZN(n1694));
  AND2_X1   g1631(.A1(358), .A2(239), .ZN(n1695));
  XNOR2_X1  g1632(.A(n1695), .B(n1694), .ZN(n1696));
  NOR2_X1   g1633(.A1(n1535), .A2(n1530), .ZN(n1697));
  NOR2_X1   g1634(.A1(n1537), .A2(n1536), .ZN(n1698));
  NOR2_X1   g1635(.A1(n1698), .A2(n1697), .ZN(n1699));
  XNOR2_X1  g1636(.A(n1699), .B(n1696), .ZN(n1700));
  AND2_X1   g1637(.A1(375), .A2(222), .ZN(n1701));
  XNOR2_X1  g1638(.A(n1701), .B(n1700), .ZN(n1702));
  NOR2_X1   g1639(.A1(n1548), .A2(n1538), .ZN(n1703));
  NOR2_X1   g1640(.A1(n1550), .A2(n1549), .ZN(n1704));
  NOR2_X1   g1641(.A1(n1704), .A2(n1703), .ZN(n1705));
  XNOR2_X1  g1642(.A(n1705), .B(n1702), .ZN(n1706));
  AND2_X1   g1643(.A1(392), .A2(205), .ZN(n1707));
  XNOR2_X1  g1644(.A(n1707), .B(n1706), .ZN(n1708));
  NOR2_X1   g1645(.A1(n1561), .A2(n1551), .ZN(n1709));
  NOR2_X1   g1646(.A1(n1563), .A2(n1562), .ZN(n1710));
  NOR2_X1   g1647(.A1(n1710), .A2(n1709), .ZN(n1711));
  XNOR2_X1  g1648(.A(n1711), .B(n1708), .ZN(n1712));
  AND2_X1   g1649(.A1(409), .A2(188), .ZN(n1713));
  XNOR2_X1  g1650(.A(n1713), .B(n1712), .ZN(n1714));
  NOR2_X1   g1651(.A1(n1574), .A2(n1564), .ZN(n1715));
  NOR2_X1   g1652(.A1(n1576), .A2(n1575), .ZN(n1716));
  NOR2_X1   g1653(.A1(n1716), .A2(n1715), .ZN(n1717));
  XNOR2_X1  g1654(.A(n1717), .B(n1714), .ZN(n1718));
  AND2_X1   g1655(.A1(426), .A2(171), .ZN(n1719));
  XNOR2_X1  g1656(.A(n1719), .B(n1718), .ZN(n1720));
  NOR2_X1   g1657(.A1(n1587), .A2(n1577), .ZN(n1721));
  NOR2_X1   g1658(.A1(n1589), .A2(n1588), .ZN(n1722));
  NOR2_X1   g1659(.A1(n1722), .A2(n1721), .ZN(n1723));
  XNOR2_X1  g1660(.A(n1723), .B(n1720), .ZN(n1724));
  AND2_X1   g1661(.A1(443), .A2(154), .ZN(n1725));
  XNOR2_X1  g1662(.A(n1725), .B(n1724), .ZN(n1726));
  NOR2_X1   g1663(.A1(n1600), .A2(n1590), .ZN(n1727));
  NOR2_X1   g1664(.A1(n1602), .A2(n1601), .ZN(n1728));
  NOR2_X1   g1665(.A1(n1728), .A2(n1727), .ZN(n1729));
  XNOR2_X1  g1666(.A(n1729), .B(n1726), .ZN(n1730));
  AND2_X1   g1667(.A1(460), .A2(137), .ZN(n1731));
  XNOR2_X1  g1668(.A(n1731), .B(n1730), .ZN(n1732));
  NOR2_X1   g1669(.A1(n1613), .A2(n1603), .ZN(n1733));
  NOR2_X1   g1670(.A1(n1615), .A2(n1614), .ZN(n1734));
  NOR2_X1   g1671(.A1(n1734), .A2(n1733), .ZN(n1735));
  XNOR2_X1  g1672(.A(n1735), .B(n1732), .ZN(n1736));
  AND2_X1   g1673(.A1(477), .A2(120), .ZN(n1737));
  XNOR2_X1  g1674(.A(n1737), .B(n1736), .ZN(n1738));
  NOR2_X1   g1675(.A1(n1626), .A2(n1616), .ZN(n1739));
  NOR2_X1   g1676(.A1(n1628), .A2(n1627), .ZN(n1740));
  NOR2_X1   g1677(.A1(n1740), .A2(n1739), .ZN(n1741));
  XNOR2_X1  g1678(.A(n1741), .B(n1738), .ZN(n1742));
  AND2_X1   g1679(.A1(494), .A2(103), .ZN(n1743));
  XNOR2_X1  g1680(.A(n1743), .B(n1742), .ZN(n1744));
  NOR2_X1   g1681(.A1(n1639), .A2(n1629), .ZN(n1745));
  NOR2_X1   g1682(.A1(n1641), .A2(n1640), .ZN(n1746));
  NOR2_X1   g1683(.A1(n1746), .A2(n1745), .ZN(n1747));
  XNOR2_X1  g1684(.A(n1747), .B(n1744), .ZN(n1748));
  AND2_X1   g1685(.A1(511), .A2(86), .ZN(n1749));
  XNOR2_X1  g1686(.A(n1749), .B(n1748), .ZN(n1750));
  NOR2_X1   g1687(.A1(n1652), .A2(n1642), .ZN(n1751));
  NOR2_X1   g1688(.A1(n1654), .A2(n1653), .ZN(n1752));
  NOR2_X1   g1689(.A1(n1752), .A2(n1751), .ZN(n1753));
  XNOR2_X1  g1690(.A(n1753), .B(n1750), .ZN(n1754));
  AND2_X1   g1691(.A1(528), .A2(69), .ZN(n1755));
  XNOR2_X1  g1692(.A(n1755), .B(n1754), .ZN(n1756));
  NOR2_X1   g1693(.A1(n1665), .A2(n1655), .ZN(n1757));
  AOI21_X1  g1694(.A(n1757), .B1(n1667), .B2(n1666), .ZN(n1758));
  XNOR2_X1  g1695(.A(n1758), .B(n1756), .ZN(n1759));
  OR2_X1    g1696(.A1(n1678), .A2(n1668), .ZN(n1760));
  OAI21_X1  g1697(.A(n1679), .B1(n1687), .B2(n1680), .ZN(n1761));
  AND2_X1   g1698(.A1(n1761), .A2(n1760), .ZN(n1762));
  XNOR2_X1  g1699(.A(n1762), .B(n1759), .ZN(6180));
  AND2_X1   g1700(.A1(358), .A2(256), .ZN(n1764));
  NOR2_X1   g1701(.A1(n1693), .A2(n1690), .ZN(n1765));
  NOR2_X1   g1702(.A1(n1695), .A2(n1694), .ZN(n1766));
  NOR2_X1   g1703(.A1(n1766), .A2(n1765), .ZN(n1767));
  XNOR2_X1  g1704(.A(n1767), .B(n1764), .ZN(n1768));
  AND2_X1   g1705(.A1(375), .A2(239), .ZN(n1769));
  XNOR2_X1  g1706(.A(n1769), .B(n1768), .ZN(n1770));
  NOR2_X1   g1707(.A1(n1699), .A2(n1696), .ZN(n1771));
  NOR2_X1   g1708(.A1(n1701), .A2(n1700), .ZN(n1772));
  NOR2_X1   g1709(.A1(n1772), .A2(n1771), .ZN(n1773));
  XNOR2_X1  g1710(.A(n1773), .B(n1770), .ZN(n1774));
  AND2_X1   g1711(.A1(392), .A2(222), .ZN(n1775));
  XNOR2_X1  g1712(.A(n1775), .B(n1774), .ZN(n1776));
  NOR2_X1   g1713(.A1(n1705), .A2(n1702), .ZN(n1777));
  NOR2_X1   g1714(.A1(n1707), .A2(n1706), .ZN(n1778));
  NOR2_X1   g1715(.A1(n1778), .A2(n1777), .ZN(n1779));
  XNOR2_X1  g1716(.A(n1779), .B(n1776), .ZN(n1780));
  AND2_X1   g1717(.A1(409), .A2(205), .ZN(n1781));
  XNOR2_X1  g1718(.A(n1781), .B(n1780), .ZN(n1782));
  NOR2_X1   g1719(.A1(n1711), .A2(n1708), .ZN(n1783));
  NOR2_X1   g1720(.A1(n1713), .A2(n1712), .ZN(n1784));
  NOR2_X1   g1721(.A1(n1784), .A2(n1783), .ZN(n1785));
  XNOR2_X1  g1722(.A(n1785), .B(n1782), .ZN(n1786));
  AND2_X1   g1723(.A1(426), .A2(188), .ZN(n1787));
  XNOR2_X1  g1724(.A(n1787), .B(n1786), .ZN(n1788));
  NOR2_X1   g1725(.A1(n1717), .A2(n1714), .ZN(n1789));
  NOR2_X1   g1726(.A1(n1719), .A2(n1718), .ZN(n1790));
  NOR2_X1   g1727(.A1(n1790), .A2(n1789), .ZN(n1791));
  XNOR2_X1  g1728(.A(n1791), .B(n1788), .ZN(n1792));
  AND2_X1   g1729(.A1(443), .A2(171), .ZN(n1793));
  XNOR2_X1  g1730(.A(n1793), .B(n1792), .ZN(n1794));
  NOR2_X1   g1731(.A1(n1723), .A2(n1720), .ZN(n1795));
  NOR2_X1   g1732(.A1(n1725), .A2(n1724), .ZN(n1796));
  NOR2_X1   g1733(.A1(n1796), .A2(n1795), .ZN(n1797));
  XNOR2_X1  g1734(.A(n1797), .B(n1794), .ZN(n1798));
  AND2_X1   g1735(.A1(460), .A2(154), .ZN(n1799));
  XNOR2_X1  g1736(.A(n1799), .B(n1798), .ZN(n1800));
  NOR2_X1   g1737(.A1(n1729), .A2(n1726), .ZN(n1801));
  NOR2_X1   g1738(.A1(n1731), .A2(n1730), .ZN(n1802));
  NOR2_X1   g1739(.A1(n1802), .A2(n1801), .ZN(n1803));
  XNOR2_X1  g1740(.A(n1803), .B(n1800), .ZN(n1804));
  AND2_X1   g1741(.A1(477), .A2(137), .ZN(n1805));
  XNOR2_X1  g1742(.A(n1805), .B(n1804), .ZN(n1806));
  NOR2_X1   g1743(.A1(n1735), .A2(n1732), .ZN(n1807));
  NOR2_X1   g1744(.A1(n1737), .A2(n1736), .ZN(n1808));
  NOR2_X1   g1745(.A1(n1808), .A2(n1807), .ZN(n1809));
  XNOR2_X1  g1746(.A(n1809), .B(n1806), .ZN(n1810));
  AND2_X1   g1747(.A1(494), .A2(120), .ZN(n1811));
  XNOR2_X1  g1748(.A(n1811), .B(n1810), .ZN(n1812));
  NOR2_X1   g1749(.A1(n1741), .A2(n1738), .ZN(n1813));
  NOR2_X1   g1750(.A1(n1743), .A2(n1742), .ZN(n1814));
  NOR2_X1   g1751(.A1(n1814), .A2(n1813), .ZN(n1815));
  XNOR2_X1  g1752(.A(n1815), .B(n1812), .ZN(n1816));
  AND2_X1   g1753(.A1(511), .A2(103), .ZN(n1817));
  XNOR2_X1  g1754(.A(n1817), .B(n1816), .ZN(n1818));
  NOR2_X1   g1755(.A1(n1747), .A2(n1744), .ZN(n1819));
  NOR2_X1   g1756(.A1(n1749), .A2(n1748), .ZN(n1820));
  NOR2_X1   g1757(.A1(n1820), .A2(n1819), .ZN(n1821));
  XOR2_X1   g1758(.A(n1821), .B(n1818), .ZN(n1822));
  NAND2_X1  g1759(.A1(528), .A2(86), .ZN(n1823));
  XNOR2_X1  g1760(.A(n1823), .B(n1822), .ZN(n1824));
  NOR2_X1   g1761(.A1(n1753), .A2(n1750), .ZN(n1825));
  NOR2_X1   g1762(.A1(n1755), .A2(n1754), .ZN(n1826));
  NOR2_X1   g1763(.A1(n1826), .A2(n1825), .ZN(n1827));
  XOR2_X1   g1764(.A(n1827), .B(n1824), .ZN(n1828));
  NOR2_X1   g1765(.A1(n1758), .A2(n1756), .ZN(n1829));
  AOI21_X1  g1766(.A(n1759), .B1(n1761), .B2(n1760), .ZN(n1830));
  OR2_X1    g1767(.A1(n1830), .A2(n1829), .ZN(n1831));
  XNOR2_X1  g1768(.A(n1831), .B(n1828), .ZN(6190));
  AND2_X1   g1769(.A1(375), .A2(256), .ZN(n1833));
  NOR2_X1   g1770(.A1(n1767), .A2(n1764), .ZN(n1834));
  NOR2_X1   g1771(.A1(n1769), .A2(n1768), .ZN(n1835));
  NOR2_X1   g1772(.A1(n1835), .A2(n1834), .ZN(n1836));
  XNOR2_X1  g1773(.A(n1836), .B(n1833), .ZN(n1837));
  AND2_X1   g1774(.A1(392), .A2(239), .ZN(n1838));
  XNOR2_X1  g1775(.A(n1838), .B(n1837), .ZN(n1839));
  NOR2_X1   g1776(.A1(n1773), .A2(n1770), .ZN(n1840));
  NOR2_X1   g1777(.A1(n1775), .A2(n1774), .ZN(n1841));
  NOR2_X1   g1778(.A1(n1841), .A2(n1840), .ZN(n1842));
  XNOR2_X1  g1779(.A(n1842), .B(n1839), .ZN(n1843));
  AND2_X1   g1780(.A1(409), .A2(222), .ZN(n1844));
  XNOR2_X1  g1781(.A(n1844), .B(n1843), .ZN(n1845));
  NOR2_X1   g1782(.A1(n1779), .A2(n1776), .ZN(n1846));
  NOR2_X1   g1783(.A1(n1781), .A2(n1780), .ZN(n1847));
  NOR2_X1   g1784(.A1(n1847), .A2(n1846), .ZN(n1848));
  XNOR2_X1  g1785(.A(n1848), .B(n1845), .ZN(n1849));
  AND2_X1   g1786(.A1(426), .A2(205), .ZN(n1850));
  XNOR2_X1  g1787(.A(n1850), .B(n1849), .ZN(n1851));
  NOR2_X1   g1788(.A1(n1785), .A2(n1782), .ZN(n1852));
  NOR2_X1   g1789(.A1(n1787), .A2(n1786), .ZN(n1853));
  NOR2_X1   g1790(.A1(n1853), .A2(n1852), .ZN(n1854));
  XNOR2_X1  g1791(.A(n1854), .B(n1851), .ZN(n1855));
  AND2_X1   g1792(.A1(443), .A2(188), .ZN(n1856));
  XNOR2_X1  g1793(.A(n1856), .B(n1855), .ZN(n1857));
  NOR2_X1   g1794(.A1(n1791), .A2(n1788), .ZN(n1858));
  NOR2_X1   g1795(.A1(n1793), .A2(n1792), .ZN(n1859));
  NOR2_X1   g1796(.A1(n1859), .A2(n1858), .ZN(n1860));
  XNOR2_X1  g1797(.A(n1860), .B(n1857), .ZN(n1861));
  AND2_X1   g1798(.A1(460), .A2(171), .ZN(n1862));
  XNOR2_X1  g1799(.A(n1862), .B(n1861), .ZN(n1863));
  NOR2_X1   g1800(.A1(n1797), .A2(n1794), .ZN(n1864));
  NOR2_X1   g1801(.A1(n1799), .A2(n1798), .ZN(n1865));
  NOR2_X1   g1802(.A1(n1865), .A2(n1864), .ZN(n1866));
  XNOR2_X1  g1803(.A(n1866), .B(n1863), .ZN(n1867));
  AND2_X1   g1804(.A1(477), .A2(154), .ZN(n1868));
  XNOR2_X1  g1805(.A(n1868), .B(n1867), .ZN(n1869));
  NOR2_X1   g1806(.A1(n1803), .A2(n1800), .ZN(n1870));
  NOR2_X1   g1807(.A1(n1805), .A2(n1804), .ZN(n1871));
  NOR2_X1   g1808(.A1(n1871), .A2(n1870), .ZN(n1872));
  XNOR2_X1  g1809(.A(n1872), .B(n1869), .ZN(n1873));
  AND2_X1   g1810(.A1(494), .A2(137), .ZN(n1874));
  XNOR2_X1  g1811(.A(n1874), .B(n1873), .ZN(n1875));
  NOR2_X1   g1812(.A1(n1809), .A2(n1806), .ZN(n1876));
  NOR2_X1   g1813(.A1(n1811), .A2(n1810), .ZN(n1877));
  NOR2_X1   g1814(.A1(n1877), .A2(n1876), .ZN(n1878));
  XNOR2_X1  g1815(.A(n1878), .B(n1875), .ZN(n1879));
  AND2_X1   g1816(.A1(511), .A2(120), .ZN(n1880));
  XNOR2_X1  g1817(.A(n1880), .B(n1879), .ZN(n1881));
  NOR2_X1   g1818(.A1(n1815), .A2(n1812), .ZN(n1882));
  NOR2_X1   g1819(.A1(n1817), .A2(n1816), .ZN(n1883));
  NOR2_X1   g1820(.A1(n1883), .A2(n1882), .ZN(n1884));
  XNOR2_X1  g1821(.A(n1884), .B(n1881), .ZN(n1885));
  AND2_X1   g1822(.A1(528), .A2(103), .ZN(n1886));
  XNOR2_X1  g1823(.A(n1886), .B(n1885), .ZN(n1887));
  NOR2_X1   g1824(.A1(n1821), .A2(n1818), .ZN(n1888));
  AOI21_X1  g1825(.A(n1888), .B1(n1823), .B2(n1822), .ZN(n1889));
  XNOR2_X1  g1826(.A(n1889), .B(n1887), .ZN(n1890));
  OR2_X1    g1827(.A1(n1827), .A2(n1824), .ZN(n1891));
  OAI21_X1  g1828(.A(n1828), .B1(n1830), .B2(n1829), .ZN(n1892));
  AND2_X1   g1829(.A1(n1892), .A2(n1891), .ZN(n1893));
  XNOR2_X1  g1830(.A(n1893), .B(n1890), .ZN(6200));
  AND2_X1   g1831(.A1(392), .A2(256), .ZN(n1895));
  NOR2_X1   g1832(.A1(n1836), .A2(n1833), .ZN(n1896));
  NOR2_X1   g1833(.A1(n1838), .A2(n1837), .ZN(n1897));
  NOR2_X1   g1834(.A1(n1897), .A2(n1896), .ZN(n1898));
  XNOR2_X1  g1835(.A(n1898), .B(n1895), .ZN(n1899));
  AND2_X1   g1836(.A1(409), .A2(239), .ZN(n1900));
  XNOR2_X1  g1837(.A(n1900), .B(n1899), .ZN(n1901));
  NOR2_X1   g1838(.A1(n1842), .A2(n1839), .ZN(n1902));
  NOR2_X1   g1839(.A1(n1844), .A2(n1843), .ZN(n1903));
  NOR2_X1   g1840(.A1(n1903), .A2(n1902), .ZN(n1904));
  XNOR2_X1  g1841(.A(n1904), .B(n1901), .ZN(n1905));
  AND2_X1   g1842(.A1(426), .A2(222), .ZN(n1906));
  XNOR2_X1  g1843(.A(n1906), .B(n1905), .ZN(n1907));
  NOR2_X1   g1844(.A1(n1848), .A2(n1845), .ZN(n1908));
  NOR2_X1   g1845(.A1(n1850), .A2(n1849), .ZN(n1909));
  NOR2_X1   g1846(.A1(n1909), .A2(n1908), .ZN(n1910));
  XNOR2_X1  g1847(.A(n1910), .B(n1907), .ZN(n1911));
  AND2_X1   g1848(.A1(443), .A2(205), .ZN(n1912));
  XNOR2_X1  g1849(.A(n1912), .B(n1911), .ZN(n1913));
  NOR2_X1   g1850(.A1(n1854), .A2(n1851), .ZN(n1914));
  NOR2_X1   g1851(.A1(n1856), .A2(n1855), .ZN(n1915));
  NOR2_X1   g1852(.A1(n1915), .A2(n1914), .ZN(n1916));
  XNOR2_X1  g1853(.A(n1916), .B(n1913), .ZN(n1917));
  AND2_X1   g1854(.A1(460), .A2(188), .ZN(n1918));
  XNOR2_X1  g1855(.A(n1918), .B(n1917), .ZN(n1919));
  NOR2_X1   g1856(.A1(n1860), .A2(n1857), .ZN(n1920));
  NOR2_X1   g1857(.A1(n1862), .A2(n1861), .ZN(n1921));
  NOR2_X1   g1858(.A1(n1921), .A2(n1920), .ZN(n1922));
  XNOR2_X1  g1859(.A(n1922), .B(n1919), .ZN(n1923));
  AND2_X1   g1860(.A1(477), .A2(171), .ZN(n1924));
  XNOR2_X1  g1861(.A(n1924), .B(n1923), .ZN(n1925));
  NOR2_X1   g1862(.A1(n1866), .A2(n1863), .ZN(n1926));
  NOR2_X1   g1863(.A1(n1868), .A2(n1867), .ZN(n1927));
  NOR2_X1   g1864(.A1(n1927), .A2(n1926), .ZN(n1928));
  XNOR2_X1  g1865(.A(n1928), .B(n1925), .ZN(n1929));
  AND2_X1   g1866(.A1(494), .A2(154), .ZN(n1930));
  XNOR2_X1  g1867(.A(n1930), .B(n1929), .ZN(n1931));
  NOR2_X1   g1868(.A1(n1872), .A2(n1869), .ZN(n1932));
  NOR2_X1   g1869(.A1(n1874), .A2(n1873), .ZN(n1933));
  NOR2_X1   g1870(.A1(n1933), .A2(n1932), .ZN(n1934));
  XNOR2_X1  g1871(.A(n1934), .B(n1931), .ZN(n1935));
  AND2_X1   g1872(.A1(511), .A2(137), .ZN(n1936));
  XNOR2_X1  g1873(.A(n1936), .B(n1935), .ZN(n1937));
  NOR2_X1   g1874(.A1(n1878), .A2(n1875), .ZN(n1938));
  NOR2_X1   g1875(.A1(n1880), .A2(n1879), .ZN(n1939));
  NOR2_X1   g1876(.A1(n1939), .A2(n1938), .ZN(n1940));
  XOR2_X1   g1877(.A(n1940), .B(n1937), .ZN(n1941));
  NAND2_X1  g1878(.A1(528), .A2(120), .ZN(n1942));
  XNOR2_X1  g1879(.A(n1942), .B(n1941), .ZN(n1943));
  NOR2_X1   g1880(.A1(n1884), .A2(n1881), .ZN(n1944));
  NOR2_X1   g1881(.A1(n1886), .A2(n1885), .ZN(n1945));
  NOR2_X1   g1882(.A1(n1945), .A2(n1944), .ZN(n1946));
  XOR2_X1   g1883(.A(n1946), .B(n1943), .ZN(n1947));
  NOR2_X1   g1884(.A1(n1889), .A2(n1887), .ZN(n1948));
  AOI21_X1  g1885(.A(n1890), .B1(n1892), .B2(n1891), .ZN(n1949));
  OR2_X1    g1886(.A1(n1949), .A2(n1948), .ZN(n1950));
  XNOR2_X1  g1887(.A(n1950), .B(n1947), .ZN(6210));
  AND2_X1   g1888(.A1(409), .A2(256), .ZN(n1952));
  NOR2_X1   g1889(.A1(n1898), .A2(n1895), .ZN(n1953));
  NOR2_X1   g1890(.A1(n1900), .A2(n1899), .ZN(n1954));
  NOR2_X1   g1891(.A1(n1954), .A2(n1953), .ZN(n1955));
  XNOR2_X1  g1892(.A(n1955), .B(n1952), .ZN(n1956));
  AND2_X1   g1893(.A1(426), .A2(239), .ZN(n1957));
  XNOR2_X1  g1894(.A(n1957), .B(n1956), .ZN(n1958));
  NOR2_X1   g1895(.A1(n1904), .A2(n1901), .ZN(n1959));
  NOR2_X1   g1896(.A1(n1906), .A2(n1905), .ZN(n1960));
  NOR2_X1   g1897(.A1(n1960), .A2(n1959), .ZN(n1961));
  XNOR2_X1  g1898(.A(n1961), .B(n1958), .ZN(n1962));
  AND2_X1   g1899(.A1(443), .A2(222), .ZN(n1963));
  XNOR2_X1  g1900(.A(n1963), .B(n1962), .ZN(n1964));
  NOR2_X1   g1901(.A1(n1910), .A2(n1907), .ZN(n1965));
  NOR2_X1   g1902(.A1(n1912), .A2(n1911), .ZN(n1966));
  NOR2_X1   g1903(.A1(n1966), .A2(n1965), .ZN(n1967));
  XNOR2_X1  g1904(.A(n1967), .B(n1964), .ZN(n1968));
  AND2_X1   g1905(.A1(460), .A2(205), .ZN(n1969));
  XNOR2_X1  g1906(.A(n1969), .B(n1968), .ZN(n1970));
  NOR2_X1   g1907(.A1(n1916), .A2(n1913), .ZN(n1971));
  NOR2_X1   g1908(.A1(n1918), .A2(n1917), .ZN(n1972));
  NOR2_X1   g1909(.A1(n1972), .A2(n1971), .ZN(n1973));
  XNOR2_X1  g1910(.A(n1973), .B(n1970), .ZN(n1974));
  AND2_X1   g1911(.A1(477), .A2(188), .ZN(n1975));
  XNOR2_X1  g1912(.A(n1975), .B(n1974), .ZN(n1976));
  NOR2_X1   g1913(.A1(n1922), .A2(n1919), .ZN(n1977));
  NOR2_X1   g1914(.A1(n1924), .A2(n1923), .ZN(n1978));
  NOR2_X1   g1915(.A1(n1978), .A2(n1977), .ZN(n1979));
  XNOR2_X1  g1916(.A(n1979), .B(n1976), .ZN(n1980));
  AND2_X1   g1917(.A1(494), .A2(171), .ZN(n1981));
  XNOR2_X1  g1918(.A(n1981), .B(n1980), .ZN(n1982));
  NOR2_X1   g1919(.A1(n1928), .A2(n1925), .ZN(n1983));
  NOR2_X1   g1920(.A1(n1930), .A2(n1929), .ZN(n1984));
  NOR2_X1   g1921(.A1(n1984), .A2(n1983), .ZN(n1985));
  XNOR2_X1  g1922(.A(n1985), .B(n1982), .ZN(n1986));
  AND2_X1   g1923(.A1(511), .A2(154), .ZN(n1987));
  XNOR2_X1  g1924(.A(n1987), .B(n1986), .ZN(n1988));
  NOR2_X1   g1925(.A1(n1934), .A2(n1931), .ZN(n1989));
  NOR2_X1   g1926(.A1(n1936), .A2(n1935), .ZN(n1990));
  NOR2_X1   g1927(.A1(n1990), .A2(n1989), .ZN(n1991));
  XNOR2_X1  g1928(.A(n1991), .B(n1988), .ZN(n1992));
  AND2_X1   g1929(.A1(528), .A2(137), .ZN(n1993));
  XNOR2_X1  g1930(.A(n1993), .B(n1992), .ZN(n1994));
  NOR2_X1   g1931(.A1(n1940), .A2(n1937), .ZN(n1995));
  AOI21_X1  g1932(.A(n1995), .B1(n1942), .B2(n1941), .ZN(n1996));
  XNOR2_X1  g1933(.A(n1996), .B(n1994), .ZN(n1997));
  OR2_X1    g1934(.A1(n1946), .A2(n1943), .ZN(n1998));
  OAI21_X1  g1935(.A(n1947), .B1(n1949), .B2(n1948), .ZN(n1999));
  AND2_X1   g1936(.A1(n1999), .A2(n1998), .ZN(n2000));
  XNOR2_X1  g1937(.A(n2000), .B(n1997), .ZN(6220));
  AND2_X1   g1938(.A1(426), .A2(256), .ZN(n2002));
  NOR2_X1   g1939(.A1(n1955), .A2(n1952), .ZN(n2003));
  NOR2_X1   g1940(.A1(n1957), .A2(n1956), .ZN(n2004));
  NOR2_X1   g1941(.A1(n2004), .A2(n2003), .ZN(n2005));
  XNOR2_X1  g1942(.A(n2005), .B(n2002), .ZN(n2006));
  AND2_X1   g1943(.A1(443), .A2(239), .ZN(n2007));
  XNOR2_X1  g1944(.A(n2007), .B(n2006), .ZN(n2008));
  NOR2_X1   g1945(.A1(n1961), .A2(n1958), .ZN(n2009));
  NOR2_X1   g1946(.A1(n1963), .A2(n1962), .ZN(n2010));
  NOR2_X1   g1947(.A1(n2010), .A2(n2009), .ZN(n2011));
  XNOR2_X1  g1948(.A(n2011), .B(n2008), .ZN(n2012));
  AND2_X1   g1949(.A1(460), .A2(222), .ZN(n2013));
  XNOR2_X1  g1950(.A(n2013), .B(n2012), .ZN(n2014));
  NOR2_X1   g1951(.A1(n1967), .A2(n1964), .ZN(n2015));
  NOR2_X1   g1952(.A1(n1969), .A2(n1968), .ZN(n2016));
  NOR2_X1   g1953(.A1(n2016), .A2(n2015), .ZN(n2017));
  XNOR2_X1  g1954(.A(n2017), .B(n2014), .ZN(n2018));
  AND2_X1   g1955(.A1(477), .A2(205), .ZN(n2019));
  XNOR2_X1  g1956(.A(n2019), .B(n2018), .ZN(n2020));
  NOR2_X1   g1957(.A1(n1973), .A2(n1970), .ZN(n2021));
  NOR2_X1   g1958(.A1(n1975), .A2(n1974), .ZN(n2022));
  NOR2_X1   g1959(.A1(n2022), .A2(n2021), .ZN(n2023));
  XNOR2_X1  g1960(.A(n2023), .B(n2020), .ZN(n2024));
  AND2_X1   g1961(.A1(494), .A2(188), .ZN(n2025));
  XNOR2_X1  g1962(.A(n2025), .B(n2024), .ZN(n2026));
  NOR2_X1   g1963(.A1(n1979), .A2(n1976), .ZN(n2027));
  NOR2_X1   g1964(.A1(n1981), .A2(n1980), .ZN(n2028));
  NOR2_X1   g1965(.A1(n2028), .A2(n2027), .ZN(n2029));
  XNOR2_X1  g1966(.A(n2029), .B(n2026), .ZN(n2030));
  AND2_X1   g1967(.A1(511), .A2(171), .ZN(n2031));
  XNOR2_X1  g1968(.A(n2031), .B(n2030), .ZN(n2032));
  NOR2_X1   g1969(.A1(n1985), .A2(n1982), .ZN(n2033));
  NOR2_X1   g1970(.A1(n1987), .A2(n1986), .ZN(n2034));
  NOR2_X1   g1971(.A1(n2034), .A2(n2033), .ZN(n2035));
  XOR2_X1   g1972(.A(n2035), .B(n2032), .ZN(n2036));
  NAND2_X1  g1973(.A1(528), .A2(154), .ZN(n2037));
  XNOR2_X1  g1974(.A(n2037), .B(n2036), .ZN(n2038));
  NOR2_X1   g1975(.A1(n1991), .A2(n1988), .ZN(n2039));
  NOR2_X1   g1976(.A1(n1993), .A2(n1992), .ZN(n2040));
  NOR2_X1   g1977(.A1(n2040), .A2(n2039), .ZN(n2041));
  XOR2_X1   g1978(.A(n2041), .B(n2038), .ZN(n2042));
  NOR2_X1   g1979(.A1(n1996), .A2(n1994), .ZN(n2043));
  AOI21_X1  g1980(.A(n1997), .B1(n1999), .B2(n1998), .ZN(n2044));
  OR2_X1    g1981(.A1(n2044), .A2(n2043), .ZN(n2045));
  XNOR2_X1  g1982(.A(n2045), .B(n2042), .ZN(6230));
  AND2_X1   g1983(.A1(443), .A2(256), .ZN(n2047));
  NOR2_X1   g1984(.A1(n2005), .A2(n2002), .ZN(n2048));
  NOR2_X1   g1985(.A1(n2007), .A2(n2006), .ZN(n2049));
  NOR2_X1   g1986(.A1(n2049), .A2(n2048), .ZN(n2050));
  XNOR2_X1  g1987(.A(n2050), .B(n2047), .ZN(n2051));
  AND2_X1   g1988(.A1(460), .A2(239), .ZN(n2052));
  XNOR2_X1  g1989(.A(n2052), .B(n2051), .ZN(n2053));
  NOR2_X1   g1990(.A1(n2011), .A2(n2008), .ZN(n2054));
  NOR2_X1   g1991(.A1(n2013), .A2(n2012), .ZN(n2055));
  NOR2_X1   g1992(.A1(n2055), .A2(n2054), .ZN(n2056));
  XNOR2_X1  g1993(.A(n2056), .B(n2053), .ZN(n2057));
  AND2_X1   g1994(.A1(477), .A2(222), .ZN(n2058));
  XNOR2_X1  g1995(.A(n2058), .B(n2057), .ZN(n2059));
  NOR2_X1   g1996(.A1(n2017), .A2(n2014), .ZN(n2060));
  NOR2_X1   g1997(.A1(n2019), .A2(n2018), .ZN(n2061));
  NOR2_X1   g1998(.A1(n2061), .A2(n2060), .ZN(n2062));
  XNOR2_X1  g1999(.A(n2062), .B(n2059), .ZN(n2063));
  AND2_X1   g2000(.A1(494), .A2(205), .ZN(n2064));
  XNOR2_X1  g2001(.A(n2064), .B(n2063), .ZN(n2065));
  NOR2_X1   g2002(.A1(n2023), .A2(n2020), .ZN(n2066));
  NOR2_X1   g2003(.A1(n2025), .A2(n2024), .ZN(n2067));
  NOR2_X1   g2004(.A1(n2067), .A2(n2066), .ZN(n2068));
  XNOR2_X1  g2005(.A(n2068), .B(n2065), .ZN(n2069));
  AND2_X1   g2006(.A1(511), .A2(188), .ZN(n2070));
  XNOR2_X1  g2007(.A(n2070), .B(n2069), .ZN(n2071));
  NOR2_X1   g2008(.A1(n2029), .A2(n2026), .ZN(n2072));
  NOR2_X1   g2009(.A1(n2031), .A2(n2030), .ZN(n2073));
  NOR2_X1   g2010(.A1(n2073), .A2(n2072), .ZN(n2074));
  XNOR2_X1  g2011(.A(n2074), .B(n2071), .ZN(n2075));
  AND2_X1   g2012(.A1(528), .A2(171), .ZN(n2076));
  XNOR2_X1  g2013(.A(n2076), .B(n2075), .ZN(n2077));
  NOR2_X1   g2014(.A1(n2035), .A2(n2032), .ZN(n2078));
  AOI21_X1  g2015(.A(n2078), .B1(n2037), .B2(n2036), .ZN(n2079));
  XNOR2_X1  g2016(.A(n2079), .B(n2077), .ZN(n2080));
  OR2_X1    g2017(.A1(n2041), .A2(n2038), .ZN(n2081));
  OAI21_X1  g2018(.A(n2042), .B1(n2044), .B2(n2043), .ZN(n2082));
  AND2_X1   g2019(.A1(n2082), .A2(n2081), .ZN(n2083));
  XNOR2_X1  g2020(.A(n2083), .B(n2080), .ZN(6240));
  AND2_X1   g2021(.A1(460), .A2(256), .ZN(n2085));
  NOR2_X1   g2022(.A1(n2050), .A2(n2047), .ZN(n2086));
  NOR2_X1   g2023(.A1(n2052), .A2(n2051), .ZN(n2087));
  NOR2_X1   g2024(.A1(n2087), .A2(n2086), .ZN(n2088));
  XNOR2_X1  g2025(.A(n2088), .B(n2085), .ZN(n2089));
  AND2_X1   g2026(.A1(477), .A2(239), .ZN(n2090));
  XNOR2_X1  g2027(.A(n2090), .B(n2089), .ZN(n2091));
  NOR2_X1   g2028(.A1(n2056), .A2(n2053), .ZN(n2092));
  NOR2_X1   g2029(.A1(n2058), .A2(n2057), .ZN(n2093));
  NOR2_X1   g2030(.A1(n2093), .A2(n2092), .ZN(n2094));
  XNOR2_X1  g2031(.A(n2094), .B(n2091), .ZN(n2095));
  AND2_X1   g2032(.A1(494), .A2(222), .ZN(n2096));
  XNOR2_X1  g2033(.A(n2096), .B(n2095), .ZN(n2097));
  NOR2_X1   g2034(.A1(n2062), .A2(n2059), .ZN(n2098));
  NOR2_X1   g2035(.A1(n2064), .A2(n2063), .ZN(n2099));
  NOR2_X1   g2036(.A1(n2099), .A2(n2098), .ZN(n2100));
  XNOR2_X1  g2037(.A(n2100), .B(n2097), .ZN(n2101));
  AND2_X1   g2038(.A1(511), .A2(205), .ZN(n2102));
  XNOR2_X1  g2039(.A(n2102), .B(n2101), .ZN(n2103));
  NOR2_X1   g2040(.A1(n2068), .A2(n2065), .ZN(n2104));
  NOR2_X1   g2041(.A1(n2070), .A2(n2069), .ZN(n2105));
  NOR2_X1   g2042(.A1(n2105), .A2(n2104), .ZN(n2106));
  XOR2_X1   g2043(.A(n2106), .B(n2103), .ZN(n2107));
  NAND2_X1  g2044(.A1(528), .A2(188), .ZN(n2108));
  XNOR2_X1  g2045(.A(n2108), .B(n2107), .ZN(n2109));
  NOR2_X1   g2046(.A1(n2074), .A2(n2071), .ZN(n2110));
  NOR2_X1   g2047(.A1(n2076), .A2(n2075), .ZN(n2111));
  NOR2_X1   g2048(.A1(n2111), .A2(n2110), .ZN(n2112));
  XOR2_X1   g2049(.A(n2112), .B(n2109), .ZN(n2113));
  NOR2_X1   g2050(.A1(n2079), .A2(n2077), .ZN(n2114));
  AOI21_X1  g2051(.A(n2080), .B1(n2082), .B2(n2081), .ZN(n2115));
  OR2_X1    g2052(.A1(n2115), .A2(n2114), .ZN(n2116));
  XNOR2_X1  g2053(.A(n2116), .B(n2113), .ZN(6250));
  AND2_X1   g2054(.A1(477), .A2(256), .ZN(n2118));
  NOR2_X1   g2055(.A1(n2088), .A2(n2085), .ZN(n2119));
  NOR2_X1   g2056(.A1(n2090), .A2(n2089), .ZN(n2120));
  NOR2_X1   g2057(.A1(n2120), .A2(n2119), .ZN(n2121));
  XNOR2_X1  g2058(.A(n2121), .B(n2118), .ZN(n2122));
  AND2_X1   g2059(.A1(494), .A2(239), .ZN(n2123));
  XNOR2_X1  g2060(.A(n2123), .B(n2122), .ZN(n2124));
  NOR2_X1   g2061(.A1(n2094), .A2(n2091), .ZN(n2125));
  NOR2_X1   g2062(.A1(n2096), .A2(n2095), .ZN(n2126));
  NOR2_X1   g2063(.A1(n2126), .A2(n2125), .ZN(n2127));
  XNOR2_X1  g2064(.A(n2127), .B(n2124), .ZN(n2128));
  AND2_X1   g2065(.A1(511), .A2(222), .ZN(n2129));
  XNOR2_X1  g2066(.A(n2129), .B(n2128), .ZN(n2130));
  NOR2_X1   g2067(.A1(n2100), .A2(n2097), .ZN(n2131));
  NOR2_X1   g2068(.A1(n2102), .A2(n2101), .ZN(n2132));
  NOR2_X1   g2069(.A1(n2132), .A2(n2131), .ZN(n2133));
  XNOR2_X1  g2070(.A(n2133), .B(n2130), .ZN(n2134));
  AND2_X1   g2071(.A1(528), .A2(205), .ZN(n2135));
  XNOR2_X1  g2072(.A(n2135), .B(n2134), .ZN(n2136));
  NOR2_X1   g2073(.A1(n2106), .A2(n2103), .ZN(n2137));
  AOI21_X1  g2074(.A(n2137), .B1(n2108), .B2(n2107), .ZN(n2138));
  XNOR2_X1  g2075(.A(n2138), .B(n2136), .ZN(n2139));
  OR2_X1    g2076(.A1(n2112), .A2(n2109), .ZN(n2140));
  OAI21_X1  g2077(.A(n2113), .B1(n2115), .B2(n2114), .ZN(n2141));
  AND2_X1   g2078(.A1(n2141), .A2(n2140), .ZN(n2142));
  XNOR2_X1  g2079(.A(n2142), .B(n2139), .ZN(6260));
  AND2_X1   g2080(.A1(494), .A2(256), .ZN(n2144));
  NOR2_X1   g2081(.A1(n2121), .A2(n2118), .ZN(n2145));
  NOR2_X1   g2082(.A1(n2123), .A2(n2122), .ZN(n2146));
  NOR2_X1   g2083(.A1(n2146), .A2(n2145), .ZN(n2147));
  XNOR2_X1  g2084(.A(n2147), .B(n2144), .ZN(n2148));
  AND2_X1   g2085(.A1(511), .A2(239), .ZN(n2149));
  XNOR2_X1  g2086(.A(n2149), .B(n2148), .ZN(n2150));
  NOR2_X1   g2087(.A1(n2127), .A2(n2124), .ZN(n2151));
  NOR2_X1   g2088(.A1(n2129), .A2(n2128), .ZN(n2152));
  NOR2_X1   g2089(.A1(n2152), .A2(n2151), .ZN(n2153));
  XOR2_X1   g2090(.A(n2153), .B(n2150), .ZN(n2154));
  NAND2_X1  g2091(.A1(528), .A2(222), .ZN(n2155));
  XNOR2_X1  g2092(.A(n2155), .B(n2154), .ZN(n2156));
  NOR2_X1   g2093(.A1(n2133), .A2(n2130), .ZN(n2157));
  NOR2_X1   g2094(.A1(n2135), .A2(n2134), .ZN(n2158));
  NOR2_X1   g2095(.A1(n2158), .A2(n2157), .ZN(n2159));
  XOR2_X1   g2096(.A(n2159), .B(n2156), .ZN(n2160));
  NOR2_X1   g2097(.A1(n2138), .A2(n2136), .ZN(n2161));
  AOI21_X1  g2098(.A(n2139), .B1(n2141), .B2(n2140), .ZN(n2162));
  OR2_X1    g2099(.A1(n2162), .A2(n2161), .ZN(n2163));
  XNOR2_X1  g2100(.A(n2163), .B(n2160), .ZN(6270));
  AND2_X1   g2101(.A1(511), .A2(256), .ZN(n2165));
  NOR2_X1   g2102(.A1(n2147), .A2(n2144), .ZN(n2166));
  NOR2_X1   g2103(.A1(n2149), .A2(n2148), .ZN(n2167));
  NOR2_X1   g2104(.A1(n2167), .A2(n2166), .ZN(n2168));
  XNOR2_X1  g2105(.A(n2168), .B(n2165), .ZN(n2169));
  AND2_X1   g2106(.A1(528), .A2(239), .ZN(n2170));
  XNOR2_X1  g2107(.A(n2170), .B(n2169), .ZN(n2171));
  NOR2_X1   g2108(.A1(n2153), .A2(n2150), .ZN(n2172));
  AOI21_X1  g2109(.A(n2172), .B1(n2155), .B2(n2154), .ZN(n2173));
  XNOR2_X1  g2110(.A(n2173), .B(n2171), .ZN(n2174));
  OR2_X1    g2111(.A1(n2159), .A2(n2156), .ZN(n2175));
  OAI21_X1  g2112(.A(n2160), .B1(n2162), .B2(n2161), .ZN(n2176));
  AND2_X1   g2113(.A1(n2176), .A2(n2175), .ZN(n2177));
  XNOR2_X1  g2114(.A(n2177), .B(n2174), .ZN(6280));
  AND2_X1   g2115(.A1(528), .A2(256), .ZN(n2179));
  NOR2_X1   g2116(.A1(n2168), .A2(n2165), .ZN(n2180));
  NOR2_X1   g2117(.A1(n2170), .A2(n2169), .ZN(n2181));
  NOR2_X1   g2118(.A1(n2181), .A2(n2180), .ZN(n2182));
  NOR2_X1   g2119(.A1(n2182), .A2(n2179), .ZN(n2183));
  INV_X1    g2120(.A(n2179), .ZN(n2184));
  XNOR2_X1  g2121(.A(n2182), .B(n2184), .ZN(n2185));
  NOR2_X1   g2122(.A1(n2173), .A2(n2171), .ZN(n2186));
  AOI21_X1  g2123(.A(n2174), .B1(n2176), .B2(n2175), .ZN(n2187));
  OR2_X1    g2124(.A1(n2187), .A2(n2186), .ZN(n2188));
  AOI21_X1  g2125(.A(n2183), .B1(n2188), .B2(n2185), .ZN(6287));
  XNOR2_X1  g2126(.A(n2188), .B(n2185), .ZN(6288));
endmodule


