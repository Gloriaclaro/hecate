// Benchmark "c432" written by ABC on Thu Dec 01 09:34:35 2022

module c432 ( 
    \1 , 4, 8, 11, 14, 17, 21, 24, 27, 30, 34, 37, 40, 43, 47, 50, 53, 56,
    60, 63, 66, 69, 73, 76, 79, 82, 86, 89, 92, 95, 99, 102, 105, 108, 112,
    115,
    223, 329, 370, 421, 430, 431, 432  );
  input  \1 , 4, 8, 11, 14, 17, 21, 24, 27, 30, 34, 37, 40, 43, 47, 50,
    53, 56, 60, 63, 66, 69, 73, 76, 79, 82, 86, 89, 92, 95, 99, 102, 105,
    108, 112, 115;
  output 223, 329, 370, 421, 430, 431, 432;
  wire n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
    n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n70, n71, n72,
    n73, n74, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
    n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n103,
    n104, n105, n109, n110, n111, n112, n113, n117, n118, n119, n123, n124,
    n125, n126, n129, n130, n131, n132, n135, n136, n137, n138, n139, n142,
    n143, n144, n145, n148, n149, n150, n151, n152, n153, n154, n158, n159,
    n160, n162, n163, n164, n165, n167, n168, n169, n170, n171, n172, n173,
    n175, n176, n177, n179, n180, n181, n182, n185, n186, n189, n190, n191,
    n194, n195, n198, n199, n200, n201, n202, n203, n204, n206, n207, n208,
    n209, n210, n213, n214, n215, n216, n217, n218, n219, n222, n223, n224,
    n225, n226, n229, n230, n231, n232, n233, n234, n237, n238, n239, n240,
    n243, n244, n245, n246, n247, n250, n251, n252, n253, n256, n257, n258,
    n259, n260, n261, n262, n264, n265, n268, n269, n272, n273, n274, n275,
    n278, n279, n282, n283, n284, n287, n288, n289, n292, n293, n294, n295,
    n298, n299, n300, n303, n304, n305, n306, n307, n308, n309, n310, n311,
    n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
    n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
    n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
    n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
    n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
    n372, n373, n374, n375, n376, n377, n378, n379, n381, n382, n383, n384,
    n385, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
    n398, n399, n400, n401, n402, n403, n404, n405, n407, n408, n409, n410,
    n411, n412, n413, n414, n415;
  INV_X1    g000(.A(108), .ZN(n43));
  NOR2_X1   g001(.A1(n43), .A2(102), .ZN(n44));
  INV_X1    g002(.A(89), .ZN(n45));
  NAND2_X1  g003(.A1(95), .A2(n45), .ZN(n46));
  INV_X1    g004(.A(76), .ZN(n47));
  NAND2_X1  g005(.A1(82), .A2(n47), .ZN(n48));
  NAND2_X1  g006(.A1(n48), .A2(n46), .ZN(n49));
  NOR2_X1   g007(.A1(n49), .A2(n44), .ZN(n50));
  INV_X1    g008(.A(\1 ), .ZN(n51));
  NAND2_X1  g009(.A1(4), .A2(n51), .ZN(n52));
  INV_X1    g010(.A(11), .ZN(n53));
  NAND2_X1  g011(.A1(17), .A2(n53), .ZN(n54));
  NAND2_X1  g012(.A1(n54), .A2(n52), .ZN(n55));
  INV_X1    g013(.A(43), .ZN(n56));
  NOR2_X1   g014(.A1(n56), .A2(37), .ZN(n57));
  INV_X1    g015(.A(30), .ZN(n58));
  NOR2_X1   g016(.A1(n58), .A2(24), .ZN(n59));
  NOR2_X1   g017(.A1(n59), .A2(n57), .ZN(n60));
  INV_X1    g018(.A(69), .ZN(n61));
  NOR2_X1   g019(.A1(n61), .A2(63), .ZN(n62));
  INV_X1    g020(.A(56), .ZN(n63));
  NOR2_X1   g021(.A1(n63), .A2(50), .ZN(n64));
  NOR2_X1   g022(.A1(n64), .A2(n62), .ZN(n65));
  NAND2_X1  g023(.A1(n65), .A2(n60), .ZN(n66));
  NOR2_X1   g024(.A1(n66), .A2(n55), .ZN(n67));
  NAND2_X1  g025(.A1(n67), .A2(n50), .ZN(223));
  INV_X1    g026(.A(95), .ZN(n70));
  NOR2_X1   g027(.A1(n70), .A2(89), .ZN(n71));
  INV_X1    g028(.A(82), .ZN(n72));
  NOR2_X1   g029(.A1(n72), .A2(76), .ZN(n73));
  NOR2_X1   g030(.A1(n73), .A2(n71), .ZN(n74));
  NOR2_X1   g031(.A1(n44), .A2(n99), .ZN(n76));
  NOR2_X1   g032(.A1(112), .A2(n43), .ZN(n77));
  INV_X1    g033(.A(n77), .ZN(n78));
  NOR2_X1   g034(.A1(n78), .A2(n76), .ZN(n79));
  INV_X1    g035(.A(n44), .ZN(n80));
  NAND2_X1  g036(.A1(n74), .A2(n80), .ZN(n81));
  INV_X1    g037(.A(4), .ZN(n82));
  NOR2_X1   g038(.A1(n82), .A2(\1 ), .ZN(n83));
  INV_X1    g039(.A(17), .ZN(n84));
  NOR2_X1   g040(.A1(n84), .A2(11), .ZN(n85));
  NOR2_X1   g041(.A1(n85), .A2(n83), .ZN(n86));
  INV_X1    g042(.A(37), .ZN(n87));
  NAND2_X1  g043(.A1(43), .A2(n87), .ZN(n88));
  INV_X1    g044(.A(24), .ZN(n89));
  NAND2_X1  g045(.A1(30), .A2(n89), .ZN(n90));
  NAND2_X1  g046(.A1(n90), .A2(n88), .ZN(n91));
  INV_X1    g047(.A(63), .ZN(n92));
  NAND2_X1  g048(.A1(69), .A2(n92), .ZN(n93));
  INV_X1    g049(.A(50), .ZN(n94));
  NAND2_X1  g050(.A1(56), .A2(n94), .ZN(n95));
  NAND2_X1  g051(.A1(n95), .A2(n93), .ZN(n96));
  NOR2_X1   g052(.A1(n96), .A2(n91), .ZN(n97));
  NAND2_X1  g053(.A1(n97), .A2(n86), .ZN(n98));
  NOR2_X1   g054(.A1(n98), .A2(n81), .ZN(n99));
  NAND2_X1  g055(.A1(n99), .A2(n46), .ZN(n100));
  NAND2_X1  g056(.A1(n46), .A2(n100), .ZN(n103));
  NOR2_X1   g057(.A1(99), .A2(n70), .ZN(n104));
  NAND2_X1  g058(.A1(n104), .A2(n103), .ZN(n105));
  NAND2_X1  g059(.A1(n48), .A2(n100), .ZN(n109));
  NOR2_X1   g060(.A1(86), .A2(n72), .ZN(n110));
  NAND2_X1  g061(.A1(n110), .A2(n109), .ZN(n111));
  NAND2_X1  g062(.A1(n111), .A2(n105), .ZN(n112));
  NOR2_X1   g063(.A1(n112), .A2(n79), .ZN(n113));
  NAND2_X1  g064(.A1(n52), .A2(n100), .ZN(n117));
  NOR2_X1   g065(.A1(8), .A2(n82), .ZN(n118));
  NAND2_X1  g066(.A1(n118), .A2(n117), .ZN(n119));
  NAND2_X1  g067(.A1(n54), .A2(n100), .ZN(n123));
  NOR2_X1   g068(.A1(21), .A2(n84), .ZN(n124));
  NAND2_X1  g069(.A1(n124), .A2(n123), .ZN(n125));
  NAND2_X1  g070(.A1(n125), .A2(n119), .ZN(n126));
  NOR2_X1   g071(.A1(n57), .A2(n99), .ZN(n129));
  NOR2_X1   g072(.A1(47), .A2(n56), .ZN(n130));
  INV_X1    g073(.A(n130), .ZN(n131));
  NOR2_X1   g074(.A1(n131), .A2(n129), .ZN(n132));
  NOR2_X1   g075(.A1(n59), .A2(n99), .ZN(n135));
  NOR2_X1   g076(.A1(34), .A2(n58), .ZN(n136));
  INV_X1    g077(.A(n136), .ZN(n137));
  NOR2_X1   g078(.A1(n137), .A2(n135), .ZN(n138));
  NOR2_X1   g079(.A1(n138), .A2(n132), .ZN(n139));
  NOR2_X1   g080(.A1(n62), .A2(n99), .ZN(n142));
  NOR2_X1   g081(.A1(73), .A2(n61), .ZN(n143));
  INV_X1    g082(.A(n143), .ZN(n144));
  NOR2_X1   g083(.A1(n144), .A2(n142), .ZN(n145));
  NOR2_X1   g084(.A1(n64), .A2(n99), .ZN(n148));
  NOR2_X1   g085(.A1(60), .A2(n63), .ZN(n149));
  INV_X1    g086(.A(n149), .ZN(n150));
  NOR2_X1   g087(.A1(n150), .A2(n148), .ZN(n151));
  NOR2_X1   g088(.A1(n151), .A2(n145), .ZN(n152));
  NAND2_X1  g089(.A1(n152), .A2(n139), .ZN(n153));
  NOR2_X1   g090(.A1(n153), .A2(n126), .ZN(n154));
  NAND2_X1  g091(.A1(n154), .A2(n113), .ZN(329));
  NOR2_X1   g092(.A1(n71), .A2(n99), .ZN(n158));
  INV_X1    g093(.A(n104), .ZN(n159));
  NOR2_X1   g094(.A1(n159), .A2(n158), .ZN(n160));
  NOR2_X1   g095(.A1(n73), .A2(n99), .ZN(n162));
  INV_X1    g096(.A(n110), .ZN(n163));
  NOR2_X1   g097(.A1(n163), .A2(n162), .ZN(n164));
  NOR2_X1   g098(.A1(n164), .A2(n160), .ZN(n165));
  NOR2_X1   g099(.A1(n79), .A2(n203), .ZN(n167));
  INV_X1    g100(.A(n76), .ZN(n168));
  NOR2_X1   g101(.A1(115), .A2(n43), .ZN(n169));
  NAND2_X1  g102(.A1(n169), .A2(n168), .ZN(n170));
  NOR2_X1   g103(.A1(n170), .A2(n167), .ZN(n171));
  INV_X1    g104(.A(n79), .ZN(n172));
  NAND2_X1  g105(.A1(n165), .A2(n172), .ZN(n173));
  NOR2_X1   g106(.A1(n83), .A2(n99), .ZN(n175));
  INV_X1    g107(.A(n118), .ZN(n176));
  NOR2_X1   g108(.A1(n176), .A2(n175), .ZN(n177));
  NOR2_X1   g109(.A1(n85), .A2(n99), .ZN(n179));
  INV_X1    g110(.A(n124), .ZN(n180));
  NOR2_X1   g111(.A1(n180), .A2(n179), .ZN(n181));
  NOR2_X1   g112(.A1(n181), .A2(n177), .ZN(n182));
  NAND2_X1  g113(.A1(n88), .A2(n100), .ZN(n185));
  NAND2_X1  g114(.A1(n130), .A2(n185), .ZN(n186));
  NAND2_X1  g115(.A1(n90), .A2(n100), .ZN(n189));
  NAND2_X1  g116(.A1(n136), .A2(n189), .ZN(n190));
  NAND2_X1  g117(.A1(n190), .A2(n186), .ZN(n191));
  NAND2_X1  g118(.A1(n93), .A2(n100), .ZN(n194));
  NAND2_X1  g119(.A1(n143), .A2(n194), .ZN(n195));
  NAND2_X1  g120(.A1(n95), .A2(n100), .ZN(n198));
  NAND2_X1  g121(.A1(n149), .A2(n198), .ZN(n199));
  NAND2_X1  g122(.A1(n199), .A2(n195), .ZN(n200));
  NOR2_X1   g123(.A1(n200), .A2(n191), .ZN(n201));
  NAND2_X1  g124(.A1(n201), .A2(n182), .ZN(n202));
  NOR2_X1   g125(.A1(n202), .A2(n173), .ZN(n203));
  NAND2_X1  g126(.A1(n203), .A2(n105), .ZN(n204));
  NAND2_X1  g127(.A1(n105), .A2(n204), .ZN(n206));
  NOR2_X1   g128(.A1(105), .A2(n70), .ZN(n207));
  NAND2_X1  g129(.A1(n207), .A2(n103), .ZN(n208));
  INV_X1    g130(.A(n208), .ZN(n209));
  NAND2_X1  g131(.A1(n209), .A2(n206), .ZN(n210));
  NAND2_X1  g132(.A1(n111), .A2(n204), .ZN(n213));
  NOR2_X1   g133(.A1(92), .A2(n72), .ZN(n214));
  NAND2_X1  g134(.A1(n214), .A2(n109), .ZN(n215));
  INV_X1    g135(.A(n215), .ZN(n216));
  NAND2_X1  g136(.A1(n216), .A2(n213), .ZN(n217));
  NAND2_X1  g137(.A1(n217), .A2(n210), .ZN(n218));
  NOR2_X1   g138(.A1(n218), .A2(n171), .ZN(n219));
  NAND2_X1  g139(.A1(n119), .A2(n204), .ZN(n222));
  NOR2_X1   g140(.A1(14), .A2(n82), .ZN(n223));
  NAND2_X1  g141(.A1(n223), .A2(n117), .ZN(n224));
  INV_X1    g142(.A(n224), .ZN(n225));
  NAND2_X1  g143(.A1(n225), .A2(n222), .ZN(n226));
  NAND2_X1  g144(.A1(n125), .A2(n204), .ZN(n229));
  NOR2_X1   g145(.A1(27), .A2(n84), .ZN(n230));
  NAND2_X1  g146(.A1(n230), .A2(n123), .ZN(n231));
  INV_X1    g147(.A(n231), .ZN(n232));
  NAND2_X1  g148(.A1(n232), .A2(n229), .ZN(n233));
  NAND2_X1  g149(.A1(n233), .A2(n226), .ZN(n234));
  NOR2_X1   g150(.A1(n132), .A2(n203), .ZN(n237));
  NOR2_X1   g151(.A1(53), .A2(n56), .ZN(n238));
  NAND2_X1  g152(.A1(n238), .A2(n185), .ZN(n239));
  NOR2_X1   g153(.A1(n239), .A2(n237), .ZN(n240));
  NOR2_X1   g154(.A1(n138), .A2(n203), .ZN(n243));
  NOR2_X1   g155(.A1(40), .A2(n58), .ZN(n244));
  NAND2_X1  g156(.A1(n244), .A2(n189), .ZN(n245));
  NOR2_X1   g157(.A1(n245), .A2(n243), .ZN(n246));
  NOR2_X1   g158(.A1(n246), .A2(n240), .ZN(n247));
  NOR2_X1   g159(.A1(n145), .A2(n203), .ZN(n250));
  NOR2_X1   g160(.A1(79), .A2(n61), .ZN(n251));
  NAND2_X1  g161(.A1(n251), .A2(n194), .ZN(n252));
  NOR2_X1   g162(.A1(n252), .A2(n250), .ZN(n253));
  NOR2_X1   g163(.A1(n151), .A2(n203), .ZN(n256));
  NOR2_X1   g164(.A1(66), .A2(n63), .ZN(n257));
  NAND2_X1  g165(.A1(n257), .A2(n198), .ZN(n258));
  NOR2_X1   g166(.A1(n258), .A2(n256), .ZN(n259));
  NOR2_X1   g167(.A1(n259), .A2(n253), .ZN(n260));
  NAND2_X1  g168(.A1(n260), .A2(n247), .ZN(n261));
  NOR2_X1   g169(.A1(n261), .A2(n234), .ZN(n262));
  NAND2_X1  g170(.A1(n262), .A2(n219), .ZN(370));
  INV_X1    g171(.A(14), .ZN(n264));
  INV_X1    g172(.A(n171), .ZN(n265));
  NOR2_X1   g173(.A1(n160), .A2(n203), .ZN(n268));
  NOR2_X1   g174(.A1(n208), .A2(n268), .ZN(n269));
  NOR2_X1   g175(.A1(n164), .A2(n203), .ZN(n272));
  NOR2_X1   g176(.A1(n215), .A2(n272), .ZN(n273));
  NOR2_X1   g177(.A1(n273), .A2(n269), .ZN(n274));
  NAND2_X1  g178(.A1(n274), .A2(n265), .ZN(n275));
  NOR2_X1   g179(.A1(n177), .A2(n203), .ZN(n278));
  NOR2_X1   g180(.A1(n224), .A2(n278), .ZN(n279));
  NOR2_X1   g181(.A1(n181), .A2(n203), .ZN(n282));
  NOR2_X1   g182(.A1(n231), .A2(n282), .ZN(n283));
  NOR2_X1   g183(.A1(n283), .A2(n279), .ZN(n284));
  NAND2_X1  g184(.A1(n186), .A2(n204), .ZN(n287));
  INV_X1    g185(.A(n239), .ZN(n288));
  NAND2_X1  g186(.A1(n288), .A2(n287), .ZN(n289));
  NAND2_X1  g187(.A1(n190), .A2(n204), .ZN(n292));
  INV_X1    g188(.A(n245), .ZN(n293));
  NAND2_X1  g189(.A1(n293), .A2(n292), .ZN(n294));
  NAND2_X1  g190(.A1(n294), .A2(n289), .ZN(n295));
  NAND2_X1  g191(.A1(n195), .A2(n204), .ZN(n298));
  INV_X1    g192(.A(n252), .ZN(n299));
  NAND2_X1  g193(.A1(n299), .A2(n298), .ZN(n300));
  NAND2_X1  g194(.A1(n199), .A2(n204), .ZN(n303));
  INV_X1    g195(.A(n258), .ZN(n304));
  NAND2_X1  g196(.A1(n304), .A2(n303), .ZN(n305));
  NAND2_X1  g197(.A1(n305), .A2(n300), .ZN(n306));
  NOR2_X1   g198(.A1(n306), .A2(n295), .ZN(n307));
  NAND2_X1  g199(.A1(n307), .A2(n284), .ZN(n308));
  NOR2_X1   g200(.A1(n308), .A2(n275), .ZN(n309));
  NOR2_X1   g201(.A1(n309), .A2(n264), .ZN(n310));
  NAND2_X1  g202(.A1(329), .A2(8), .ZN(n311));
  NOR2_X1   g203(.A1(n99), .A2(n51), .ZN(n312));
  NOR2_X1   g204(.A1(n312), .A2(n82), .ZN(n313));
  NAND2_X1  g205(.A1(n313), .A2(n311), .ZN(n314));
  NOR2_X1   g206(.A1(n314), .A2(n310), .ZN(n315));
  INV_X1    g207(.A(66), .ZN(n316));
  NOR2_X1   g208(.A1(n309), .A2(n316), .ZN(n317));
  NAND2_X1  g209(.A1(329), .A2(60), .ZN(n318));
  NOR2_X1   g210(.A1(n99), .A2(n94), .ZN(n319));
  NOR2_X1   g211(.A1(n319), .A2(n63), .ZN(n320));
  NAND2_X1  g212(.A1(n320), .A2(n318), .ZN(n321));
  NOR2_X1   g213(.A1(n321), .A2(n317), .ZN(n322));
  INV_X1    g214(.A(53), .ZN(n323));
  NOR2_X1   g215(.A1(n309), .A2(n323), .ZN(n324));
  NAND2_X1  g216(.A1(329), .A2(47), .ZN(n325));
  NOR2_X1   g217(.A1(n99), .A2(n87), .ZN(n326));
  NOR2_X1   g218(.A1(n326), .A2(n56), .ZN(n327));
  NAND2_X1  g219(.A1(n327), .A2(n325), .ZN(n328));
  NOR2_X1   g220(.A1(n328), .A2(n324), .ZN(n329));
  NOR2_X1   g221(.A1(n329), .A2(n322), .ZN(n330));
  INV_X1    g222(.A(92), .ZN(n331));
  NOR2_X1   g223(.A1(n309), .A2(n331), .ZN(n332));
  NAND2_X1  g224(.A1(329), .A2(86), .ZN(n333));
  NOR2_X1   g225(.A1(n99), .A2(n47), .ZN(n334));
  NOR2_X1   g226(.A1(n334), .A2(n72), .ZN(n335));
  NAND2_X1  g227(.A1(n335), .A2(n333), .ZN(n336));
  NOR2_X1   g228(.A1(n336), .A2(n332), .ZN(n337));
  INV_X1    g229(.A(79), .ZN(n338));
  NOR2_X1   g230(.A1(n309), .A2(n338), .ZN(n339));
  NAND2_X1  g231(.A1(329), .A2(73), .ZN(n340));
  NOR2_X1   g232(.A1(n99), .A2(n92), .ZN(n341));
  NOR2_X1   g233(.A1(n341), .A2(n61), .ZN(n342));
  NAND2_X1  g234(.A1(n342), .A2(n340), .ZN(n343));
  NOR2_X1   g235(.A1(n343), .A2(n339), .ZN(n344));
  NOR2_X1   g236(.A1(n344), .A2(n337), .ZN(n345));
  NAND2_X1  g237(.A1(n345), .A2(n330), .ZN(n346));
  INV_X1    g238(.A(27), .ZN(n347));
  NOR2_X1   g239(.A1(n309), .A2(n347), .ZN(n348));
  NAND2_X1  g240(.A1(329), .A2(21), .ZN(n349));
  NOR2_X1   g241(.A1(n99), .A2(n53), .ZN(n350));
  NOR2_X1   g242(.A1(n350), .A2(n84), .ZN(n351));
  NAND2_X1  g243(.A1(n351), .A2(n349), .ZN(n352));
  NOR2_X1   g244(.A1(n352), .A2(n348), .ZN(n353));
  INV_X1    g245(.A(40), .ZN(n354));
  NOR2_X1   g246(.A1(n309), .A2(n354), .ZN(n355));
  NAND2_X1  g247(.A1(329), .A2(34), .ZN(n356));
  NOR2_X1   g248(.A1(n99), .A2(n89), .ZN(n357));
  NOR2_X1   g249(.A1(n357), .A2(n58), .ZN(n358));
  NAND2_X1  g250(.A1(n358), .A2(n356), .ZN(n359));
  NOR2_X1   g251(.A1(n359), .A2(n355), .ZN(n360));
  NOR2_X1   g252(.A1(n360), .A2(n353), .ZN(n361));
  INV_X1    g253(.A(115), .ZN(n362));
  NOR2_X1   g254(.A1(n309), .A2(n362), .ZN(n363));
  NAND2_X1  g255(.A1(329), .A2(112), .ZN(n364));
  INV_X1    g256(.A(102), .ZN(n365));
  NOR2_X1   g257(.A1(n99), .A2(n365), .ZN(n366));
  NOR2_X1   g258(.A1(n366), .A2(n43), .ZN(n367));
  NAND2_X1  g259(.A1(n367), .A2(n364), .ZN(n368));
  NOR2_X1   g260(.A1(n368), .A2(n363), .ZN(n369));
  INV_X1    g261(.A(105), .ZN(n370));
  NOR2_X1   g262(.A1(n309), .A2(n370), .ZN(n371));
  NAND2_X1  g263(.A1(329), .A2(99), .ZN(n372));
  NOR2_X1   g264(.A1(n99), .A2(n45), .ZN(n373));
  NOR2_X1   g265(.A1(n373), .A2(n70), .ZN(n374));
  NAND2_X1  g266(.A1(n374), .A2(n372), .ZN(n375));
  NOR2_X1   g267(.A1(n375), .A2(n371), .ZN(n376));
  NOR2_X1   g268(.A1(n376), .A2(n369), .ZN(n377));
  NAND2_X1  g269(.A1(n377), .A2(n361), .ZN(n378));
  NOR2_X1   g270(.A1(n378), .A2(n346), .ZN(n379));
  NOR2_X1   g271(.A1(n379), .A2(n315), .ZN(421));
  NAND2_X1  g272(.A1(370), .A2(53), .ZN(n381));
  INV_X1    g273(.A(n328), .ZN(n382));
  NAND2_X1  g274(.A1(n382), .A2(n381), .ZN(n383));
  NOR2_X1   g275(.A1(n360), .A2(n383), .ZN(n384));
  NOR2_X1   g276(.A1(n384), .A2(n322), .ZN(n385));
  NAND2_X1  g277(.A1(n385), .A2(n361), .ZN(430));
  NOR2_X1   g278(.A1(n360), .A2(n329), .ZN(n387));
  NAND2_X1  g279(.A1(370), .A2(79), .ZN(n388));
  INV_X1    g280(.A(n343), .ZN(n389));
  NAND2_X1  g281(.A1(n389), .A2(n388), .ZN(n390));
  NOR2_X1   g282(.A1(n390), .A2(n322), .ZN(n391));
  NAND2_X1  g283(.A1(n391), .A2(n387), .ZN(n392));
  NAND2_X1  g284(.A1(370), .A2(27), .ZN(n393));
  INV_X1    g285(.A(n352), .ZN(n394));
  NAND2_X1  g286(.A1(n394), .A2(n393), .ZN(n395));
  NAND2_X1  g287(.A1(370), .A2(40), .ZN(n396));
  INV_X1    g288(.A(n359), .ZN(n397));
  NAND2_X1  g289(.A1(n397), .A2(n396), .ZN(n398));
  NAND2_X1  g290(.A1(n398), .A2(n395), .ZN(n399));
  NAND2_X1  g291(.A1(370), .A2(66), .ZN(n400));
  INV_X1    g292(.A(n321), .ZN(n401));
  NAND2_X1  g293(.A1(n401), .A2(n400), .ZN(n402));
  NAND2_X1  g294(.A1(n337), .A2(n402), .ZN(n403));
  NOR2_X1   g295(.A1(n403), .A2(n329), .ZN(n404));
  NOR2_X1   g296(.A1(n404), .A2(n399), .ZN(n405));
  NAND2_X1  g297(.A1(n405), .A2(n392), .ZN(431));
  NAND2_X1  g298(.A1(n398), .A2(n383), .ZN(n407));
  NAND2_X1  g299(.A1(370), .A2(92), .ZN(n408));
  INV_X1    g300(.A(n336), .ZN(n409));
  NAND2_X1  g301(.A1(n409), .A2(n408), .ZN(n410));
  NAND2_X1  g302(.A1(n376), .A2(n410), .ZN(n411));
  NOR2_X1   g303(.A1(n411), .A2(n407), .ZN(n412));
  NAND2_X1  g304(.A1(n398), .A2(n329), .ZN(n413));
  NAND2_X1  g305(.A1(n413), .A2(n395), .ZN(n414));
  NOR2_X1   g306(.A1(n414), .A2(n412), .ZN(n415));
  NAND2_X1  g307(.A1(n415), .A2(n392), .ZN(432));
endmodule


