// Benchmark "c3540" written by ABC on Wed Oct 05 14:32:33 2022

module c3540 ( 
    \1 , 13, 20, 33, 41, 45, 50, 58, 68, 77, 87, 97, 107, 116, 124, 125,
    128, 132, 137, 143, 150, 159, 169, 179, 190, 200, 213, 222, 223, 226,
    232, 238, 244, 250, 257, 264, 270, 274, 283, 294, 303, 311, 317, 322,
    326, 329, 330, 343, 349, 350,
    1713, 1947, 3195, 3833, 3987, 4028, 4145, 4589, 4667, 4815, 4944, 5002,
    5045, 5047, 5078, 5102, 5120, 5121, 5192, 5231, 5360, 5361  );
  input  \1 , 13, 20, 33, 41, 45, 50, 58, 68, 77, 87, 97, 107, 116, 124,
    125, 128, 132, 137, 143, 150, 159, 169, 179, 190, 200, 213, 222, 223,
    226, 232, 238, 244, 250, 257, 264, 270, 274, 283, 294, 303, 311, 317,
    322, 326, 329, 330, 343, 349, 350;
  output 1713, 1947, 3195, 3833, 3987, 4028, 4145, 4589, 4667, 4815, 4944,
    5002, 5045, 5047, 5078, 5102, 5120, 5121, 5192, 5231, 5360, 5361;
  wire n73, n74, n75, n76, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
    n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n101, n102,
    n103, n104, n105, n106, n108, n109, n110, n111, n112, n113, n115, n116,
    n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
    n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
    n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
    n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
    n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
    n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
    n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
    n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
    n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
    n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
    n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
    n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
    n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
    n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
    n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
    n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
    n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
    n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
    n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
    n347, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
    n360, n361, n362, n364, n365, n366, n367, n368, n369, n370, n371, n372,
    n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
    n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
    n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
    n409, n410, n411, n412, n414, n415, n416, n417, n418, n419, n420, n421,
    n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
    n434, n435, n436, n437, n438, n439, n441, n442, n443, n444, n445, n446,
    n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
    n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n470, n471,
    n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
    n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
    n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
    n508, n509, n510, n511, n513, n514, n515, n516, n517, n518, n519, n520,
    n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
    n533, n534, n535, n537, n538, n539, n540, n541, n542, n543, n544, n545,
    n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n558,
    n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
    n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
    n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
    n595, n596, n597, n599, n600, n601, n602, n603, n604, n605, n606, n607,
    n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
    n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
    n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
    n644, n645, n646, n648, n649, n650, n651, n652, n653, n654, n655, n656,
    n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
    n669, n671, n672, n674, n675, n677, n678, n679, n680, n681, n682, n683,
    n684, n685, n686, n687, n688, n689, n690, n691, n693, n694;
  NOR4_X1   g000(.A1(68), .A2(58), .A3(50), .A4(77), .ZN(1713));
  INV_X1    g001(.A(87), .ZN(n73));
  INV_X1    g002(.A(97), .ZN(n74));
  INV_X1    g003(.A(107), .ZN(n75));
  AOI21_X1  g004(.A(n73), .B1(n75), .B2(n74), .ZN(n76));
  INV_X1    g005(.A(n76), .ZN(1947));
  AND3_X1   g006(.A1(20), .A2(13), .A3(\1 ), .ZN(n78));
  INV_X1    g007(.A(\1 ), .ZN(n79));
  INV_X1    g008(.A(20), .ZN(n80));
  NOR3_X1   g009(.A1(n80), .A2(13), .A3(n79), .ZN(n81));
  INV_X1    g010(.A(50), .ZN(n82));
  INV_X1    g011(.A(68), .ZN(n83));
  INV_X1    g012(.A(226), .ZN(n84));
  INV_X1    g013(.A(238), .ZN(n85));
  AOI22_X1  g014(.A1(232), .A2(58), .B1(116), .B2(270), .ZN(n86));
  OAI221_X1 g015(.A(n86), .B1(n84), .B2(n82), .C1(n83), .C2(n85), .ZN(n87));
  INV_X1    g016(.A(77), .ZN(n88));
  INV_X1    g017(.A(244), .ZN(n89));
  INV_X1    g018(.A(257), .ZN(n90));
  AOI22_X1  g019(.A1(250), .A2(87), .B1(107), .B2(264), .ZN(n91));
  OAI221_X1 g020(.A(n91), .B1(n89), .B2(n88), .C1(n74), .C2(n90), .ZN(n92));
  NOR2_X1   g021(.A1(n92), .A2(n87), .ZN(n93));
  NOR3_X1   g022(.A1(n81), .A2(n78), .A3(n93), .ZN(n94));
  INV_X1    g023(.A(58), .ZN(n95));
  AOI21_X1  g024(.A(n82), .B1(n83), .B2(n95), .ZN(n96));
  INV_X1    g025(.A(250), .ZN(n97));
  INV_X1    g026(.A(264), .ZN(n98));
  AOI21_X1  g027(.A(n97), .B1(n98), .B2(n90), .ZN(n99));
  AOI221_X1 g028(.A(n94), .B1(n81), .B2(n99), .C1(n78), .C2(n96), .ZN(3195));
  XNOR2_X1  g029(.A(270), .B(264), .ZN(n101));
  XNOR2_X1  g030(.A(257), .B(250), .ZN(n102));
  XNOR2_X1  g031(.A(n102), .B(n101), .ZN(n103));
  XNOR2_X1  g032(.A(244), .B(238), .ZN(n104));
  XNOR2_X1  g033(.A(232), .B(226), .ZN(n105));
  XNOR2_X1  g034(.A(n105), .B(n104), .ZN(n106));
  XNOR2_X1  g035(.A(n106), .B(n103), .ZN(3833));
  XNOR2_X1  g036(.A(116), .B(107), .ZN(n108));
  XNOR2_X1  g037(.A(97), .B(87), .ZN(n109));
  XNOR2_X1  g038(.A(n109), .B(n108), .ZN(n110));
  XNOR2_X1  g039(.A(77), .B(68), .ZN(n111));
  XOR2_X1   g040(.A(58), .B(50), .ZN(n112));
  XNOR2_X1  g041(.A(n112), .B(n111), .ZN(n113));
  XOR2_X1   g042(.A(n113), .B(n110), .ZN(3987));
  NAND2_X1  g043(.A1(13), .A2(\1 ), .ZN(n115));
  NAND3_X1  g044(.A1(33), .A2(20), .A3(\1 ), .ZN(n116));
  AND2_X1   g045(.A1(n116), .A2(n115), .ZN(n117));
  OR3_X1    g046(.A1(107), .A2(97), .A3(87), .ZN(n118));
  NAND2_X1  g047(.A1(n118), .A2(20), .ZN(n119));
  INV_X1    g048(.A(33), .ZN(n120));
  NAND3_X1  g049(.A1(68), .A2(n120), .A3(n80), .ZN(n121));
  NAND3_X1  g050(.A1(97), .A2(33), .A3(n80), .ZN(n122));
  AND3_X1   g051(.A1(n122), .A2(n121), .A3(n119), .ZN(n123));
  NAND3_X1  g052(.A1(20), .A2(13), .A3(n79), .ZN(n124));
  NAND2_X1  g053(.A1(33), .A2(n79), .ZN(n125));
  NAND4_X1  g054(.A1(n124), .A2(n117), .A3(87), .A4(n125), .ZN(n126));
  OAI221_X1 g055(.A(n126), .B1(n123), .B2(n117), .C1(87), .C2(n124), .ZN(n127));
  AND2_X1   g056(.A1(13), .A2(\1 ), .ZN(n128));
  NAND2_X1  g057(.A1(41), .A2(33), .ZN(n129));
  NAND2_X1  g058(.A1(n129), .A2(n128), .ZN(n130));
  NAND3_X1  g059(.A1(349), .A2(244), .A3(n120), .ZN(n131));
  NOR2_X1   g060(.A1(349), .A2(33), .ZN(n132));
  AOI22_X1  g061(.A1(238), .A2(n132), .B1(116), .B2(33), .ZN(n133));
  AOI21_X1  g062(.A(n130), .B1(n133), .B2(n131), .ZN(n134));
  AOI221_X1 g063(.A(n97), .B1(45), .B2(n79), .C1(n129), .C2(n128), .ZN(n135));
  INV_X1    g064(.A(45), .ZN(n136));
  AND2_X1   g065(.A1(41), .A2(33), .ZN(n137));
  OAI21_X1  g066(.A(274), .B1(n137), .B2(n115), .ZN(n138));
  NOR3_X1   g067(.A1(n138), .A2(n136), .A3(\1 ), .ZN(n139));
  OR3_X1    g068(.A1(n139), .A2(n135), .A3(n134), .ZN(n140));
  NAND3_X1  g069(.A1(n140), .A2(n127), .A3(169), .ZN(n141));
  NOR3_X1   g070(.A1(n139), .A2(n135), .A3(n134), .ZN(n142));
  NAND3_X1  g071(.A1(n142), .A2(n127), .A3(179), .ZN(n143));
  INV_X1    g072(.A(190), .ZN(n144));
  NOR3_X1   g073(.A1(n140), .A2(n127), .A3(n144), .ZN(n145));
  INV_X1    g074(.A(200), .ZN(n146));
  NAND2_X1  g075(.A1(n116), .A2(n115), .ZN(n147));
  NAND3_X1  g076(.A1(n122), .A2(n121), .A3(n119), .ZN(n148));
  INV_X1    g077(.A(13), .ZN(n149));
  NOR3_X1   g078(.A1(n80), .A2(n149), .A3(\1 ), .ZN(n150));
  NOR2_X1   g079(.A1(n120), .A2(\1 ), .ZN(n151));
  NOR4_X1   g080(.A1(n150), .A2(n147), .A3(n73), .A4(n151), .ZN(n152));
  AOI221_X1 g081(.A(n152), .B1(n148), .B2(n147), .C1(n73), .C2(n150), .ZN(n153));
  OAI21_X1  g082(.A(n153), .B1(n142), .B2(n146), .ZN(n154));
  OAI211_X1 g083(.A(n143), .B(n141), .C1(n145), .C2(n154), .ZN(n155));
  INV_X1    g084(.A(169), .ZN(n156));
  NAND2_X1  g085(.A1(33), .A2(n80), .ZN(n157));
  XOR2_X1   g086(.A(107), .B(97), .ZN(n158));
  NAND3_X1  g087(.A1(77), .A2(n120), .A3(n80), .ZN(n159));
  OAI221_X1 g088(.A(n159), .B1(n157), .B2(n75), .C1(n80), .C2(n158), .ZN(n160));
  NOR4_X1   g089(.A1(n150), .A2(n147), .A3(n74), .A4(n151), .ZN(n161));
  AOI221_X1 g090(.A(n161), .B1(n150), .B2(n74), .C1(n147), .C2(n160), .ZN(n162));
  NOR2_X1   g091(.A1(n137), .A2(n115), .ZN(n163));
  INV_X1    g092(.A(349), .ZN(n164));
  NOR3_X1   g093(.A1(n164), .A2(n97), .A3(33), .ZN(n165));
  INV_X1    g094(.A(283), .ZN(n166));
  OR2_X1    g095(.A1(349), .A2(33), .ZN(n167));
  OAI22_X1  g096(.A1(n166), .A2(n120), .B1(n89), .B2(n167), .ZN(n168));
  OAI21_X1  g097(.A(n163), .B1(n168), .B2(n165), .ZN(n169));
  INV_X1    g098(.A(41), .ZN(n170));
  NAND3_X1  g099(.A1(45), .A2(n170), .A3(n79), .ZN(n171));
  OR2_X1    g100(.A1(n171), .A2(n138), .ZN(n172));
  NAND3_X1  g101(.A1(n171), .A2(n130), .A3(257), .ZN(n173));
  AND3_X1   g102(.A1(n173), .A2(n172), .A3(n169), .ZN(n174));
  OR3_X1    g103(.A1(n174), .A2(n162), .A3(n156), .ZN(n175));
  NAND4_X1  g104(.A1(n172), .A2(n169), .A3(179), .A4(n173), .ZN(n176));
  OR2_X1    g105(.A1(n176), .A2(n162), .ZN(n177));
  AND3_X1   g106(.A1(n174), .A2(n162), .A3(190), .ZN(n178));
  OAI21_X1  g107(.A(n162), .B1(n174), .B2(n146), .ZN(n179));
  OAI211_X1 g108(.A(n177), .B(n175), .C1(n178), .C2(n179), .ZN(n180));
  NOR2_X1   g109(.A1(n180), .A2(n155), .ZN(n181));
  INV_X1    g110(.A(116), .ZN(n182));
  NAND3_X1  g111(.A1(97), .A2(n120), .A3(n80), .ZN(n183));
  OAI221_X1 g112(.A(n183), .B1(n166), .B2(n157), .C1(n182), .C2(n80), .ZN(n184));
  NOR4_X1   g113(.A1(n150), .A2(n147), .A3(n182), .A4(n151), .ZN(n185));
  AOI221_X1 g114(.A(n185), .B1(n150), .B2(n182), .C1(n147), .C2(n184), .ZN(n186));
  NOR3_X1   g115(.A1(n164), .A2(n98), .A3(33), .ZN(n187));
  INV_X1    g116(.A(303), .ZN(n188));
  OAI22_X1  g117(.A1(n188), .A2(n120), .B1(n90), .B2(n167), .ZN(n189));
  OAI21_X1  g118(.A(n163), .B1(n189), .B2(n187), .ZN(n190));
  NAND3_X1  g119(.A1(n171), .A2(n130), .A3(270), .ZN(n191));
  AND3_X1   g120(.A1(n191), .A2(n190), .A3(n172), .ZN(n192));
  NOR3_X1   g121(.A1(n192), .A2(n186), .A3(n156), .ZN(n193));
  INV_X1    g122(.A(179), .ZN(n194));
  NAND3_X1  g123(.A1(n191), .A2(n190), .A3(n172), .ZN(n195));
  NOR3_X1   g124(.A1(n195), .A2(n186), .A3(n194), .ZN(n196));
  OR2_X1    g125(.A1(n196), .A2(n193), .ZN(n197));
  NAND3_X1  g126(.A1(n192), .A2(n186), .A3(190), .ZN(n198));
  NAND3_X1  g127(.A1(n195), .A2(n186), .A3(200), .ZN(n199));
  AND3_X1   g128(.A1(n199), .A2(n198), .A3(n186), .ZN(n200));
  NOR2_X1   g129(.A1(n120), .A2(20), .ZN(n201));
  NOR3_X1   g130(.A1(n73), .A2(33), .A3(20), .ZN(n202));
  AOI221_X1 g131(.A(n202), .B1(116), .B2(n201), .C1(n75), .C2(20), .ZN(n203));
  NAND4_X1  g132(.A1(n124), .A2(n117), .A3(107), .A4(n125), .ZN(n204));
  OAI221_X1 g133(.A(n204), .B1(n124), .B2(107), .C1(n117), .C2(n203), .ZN(n205));
  NOR3_X1   g134(.A1(n164), .A2(n90), .A3(33), .ZN(n206));
  INV_X1    g135(.A(294), .ZN(n207));
  OAI22_X1  g136(.A1(n207), .A2(n120), .B1(n97), .B2(n167), .ZN(n208));
  OAI21_X1  g137(.A(n163), .B1(n208), .B2(n206), .ZN(n209));
  NAND3_X1  g138(.A1(n171), .A2(n130), .A3(264), .ZN(n210));
  NAND3_X1  g139(.A1(n210), .A2(n209), .A3(n172), .ZN(n211));
  NAND3_X1  g140(.A1(n211), .A2(n205), .A3(169), .ZN(n212));
  AND3_X1   g141(.A1(n210), .A2(n209), .A3(n172), .ZN(n213));
  NAND3_X1  g142(.A1(n213), .A2(n205), .A3(179), .ZN(n214));
  NOR3_X1   g143(.A1(n211), .A2(n205), .A3(n144), .ZN(n215));
  NAND3_X1  g144(.A1(87), .A2(n120), .A3(n80), .ZN(n216));
  OAI221_X1 g145(.A(n216), .B1(n182), .B2(n157), .C1(107), .C2(n80), .ZN(n217));
  NOR4_X1   g146(.A1(n150), .A2(n147), .A3(n75), .A4(n151), .ZN(n218));
  AOI221_X1 g147(.A(n218), .B1(n150), .B2(n75), .C1(n147), .C2(n217), .ZN(n219));
  OAI21_X1  g148(.A(n219), .B1(n213), .B2(n146), .ZN(n220));
  OAI211_X1 g149(.A(n214), .B(n212), .C1(n215), .C2(n220), .ZN(n221));
  NOR3_X1   g150(.A1(n221), .A2(n200), .A3(n197), .ZN(n222));
  NAND2_X1  g151(.A1(n222), .A2(n181), .ZN(n223));
  NOR3_X1   g152(.A1(68), .A2(58), .A3(50), .ZN(n224));
  NAND3_X1  g153(.A1(150), .A2(n120), .A3(n80), .ZN(n225));
  OAI221_X1 g154(.A(n225), .B1(n224), .B2(n80), .C1(n95), .C2(n157), .ZN(n226));
  NOR2_X1   g155(.A1(n80), .A2(\1 ), .ZN(n227));
  NOR4_X1   g156(.A1(n227), .A2(n147), .A3(n82), .A4(n150), .ZN(n228));
  AOI221_X1 g157(.A(n228), .B1(n150), .B2(n82), .C1(n147), .C2(n226), .ZN(n229));
  NAND3_X1  g158(.A1(349), .A2(223), .A3(n120), .ZN(n230));
  AOI22_X1  g159(.A1(222), .A2(n132), .B1(77), .B2(33), .ZN(n231));
  AOI21_X1  g160(.A(n130), .B1(n231), .B2(n230), .ZN(n232));
  OR2_X1    g161(.A1(45), .A2(41), .ZN(n233));
  NAND2_X1  g162(.A1(n233), .A2(n79), .ZN(n234));
  NOR2_X1   g163(.A1(45), .A2(41), .ZN(n235));
  OAI221_X1 g164(.A(226), .B1(n115), .B2(n137), .C1(\1 ), .C2(n235), .ZN(n236));
  OAI21_X1  g165(.A(n236), .B1(n234), .B2(n138), .ZN(n237));
  NOR2_X1   g166(.A1(n237), .A2(n232), .ZN(n238));
  NOR3_X1   g167(.A1(n238), .A2(n229), .A3(n156), .ZN(n239));
  NOR4_X1   g168(.A1(n232), .A2(n229), .A3(n194), .A4(n237), .ZN(n240));
  NOR2_X1   g169(.A1(n240), .A2(n239), .ZN(n241));
  OR3_X1    g170(.A1(n237), .A2(n232), .A3(n144), .ZN(n242));
  OAI211_X1 g171(.A(n229), .B(n242), .C1(n238), .C2(n146), .ZN(n243));
  NAND2_X1  g172(.A1(n243), .A2(n241), .ZN(n244));
  XOR2_X1   g173(.A(68), .B(58), .ZN(n245));
  NOR2_X1   g174(.A1(n245), .A2(n80), .ZN(n246));
  INV_X1    g175(.A(159), .ZN(n247));
  NOR3_X1   g176(.A1(n247), .A2(33), .A3(20), .ZN(n248));
  NOR3_X1   g177(.A1(n83), .A2(n120), .A3(20), .ZN(n249));
  NOR3_X1   g178(.A1(n249), .A2(n248), .A3(n246), .ZN(n250));
  NAND2_X1  g179(.A1(20), .A2(n79), .ZN(n251));
  NAND4_X1  g180(.A1(n251), .A2(n117), .A3(58), .A4(n124), .ZN(n252));
  OAI221_X1 g181(.A(n252), .B1(n124), .B2(58), .C1(n117), .C2(n250), .ZN(n253));
  NOR3_X1   g182(.A1(n164), .A2(n84), .A3(33), .ZN(n254));
  INV_X1    g183(.A(223), .ZN(n255));
  OAI22_X1  g184(.A1(n255), .A2(n167), .B1(n73), .B2(n120), .ZN(n256));
  OAI21_X1  g185(.A(n163), .B1(n256), .B2(n254), .ZN(n257));
  INV_X1    g186(.A(274), .ZN(n258));
  AOI21_X1  g187(.A(n258), .B1(n129), .B2(n128), .ZN(n259));
  NOR2_X1   g188(.A1(n235), .A2(\1 ), .ZN(n260));
  INV_X1    g189(.A(232), .ZN(n261));
  AOI221_X1 g190(.A(n261), .B1(n128), .B2(n129), .C1(n79), .C2(n233), .ZN(n262));
  AOI21_X1  g191(.A(n262), .B1(n260), .B2(n259), .ZN(n263));
  AOI21_X1  g192(.A(n156), .B1(n263), .B2(n257), .ZN(n264));
  NAND3_X1  g193(.A1(349), .A2(226), .A3(n120), .ZN(n265));
  AOI22_X1  g194(.A1(223), .A2(n132), .B1(87), .B2(33), .ZN(n266));
  AOI21_X1  g195(.A(n130), .B1(n266), .B2(n265), .ZN(n267));
  OAI221_X1 g196(.A(232), .B1(n115), .B2(n137), .C1(\1 ), .C2(n235), .ZN(n268));
  OAI21_X1  g197(.A(n268), .B1(n234), .B2(n138), .ZN(n269));
  NOR3_X1   g198(.A1(n269), .A2(n267), .A3(n194), .ZN(n270));
  OAI21_X1  g199(.A(n253), .B1(n270), .B2(n264), .ZN(n271));
  OR3_X1    g200(.A1(n249), .A2(n248), .A3(n246), .ZN(n272));
  NOR4_X1   g201(.A1(n227), .A2(n147), .A3(n95), .A4(n150), .ZN(n273));
  AOI221_X1 g202(.A(n273), .B1(n150), .B2(n95), .C1(n147), .C2(n272), .ZN(n274));
  NOR2_X1   g203(.A1(n269), .A2(n267), .ZN(n275));
  AND3_X1   g204(.A1(n275), .A2(n274), .A3(190), .ZN(n276));
  OAI21_X1  g205(.A(n274), .B1(n275), .B2(n146), .ZN(n277));
  OAI21_X1  g206(.A(n271), .B1(n277), .B2(n276), .ZN(n278));
  NAND3_X1  g207(.A1(58), .A2(n120), .A3(n80), .ZN(n279));
  OAI221_X1 g208(.A(n279), .B1(n73), .B2(n157), .C1(n88), .C2(n80), .ZN(n280));
  NOR4_X1   g209(.A1(n227), .A2(n147), .A3(n88), .A4(n150), .ZN(n281));
  AOI221_X1 g210(.A(n281), .B1(n150), .B2(n88), .C1(n147), .C2(n280), .ZN(n282));
  NAND3_X1  g211(.A1(349), .A2(238), .A3(n120), .ZN(n283));
  AOI22_X1  g212(.A1(232), .A2(n132), .B1(107), .B2(33), .ZN(n284));
  AOI21_X1  g213(.A(n130), .B1(n284), .B2(n283), .ZN(n285));
  OAI221_X1 g214(.A(244), .B1(n115), .B2(n137), .C1(\1 ), .C2(n235), .ZN(n286));
  OAI21_X1  g215(.A(n286), .B1(n234), .B2(n138), .ZN(n287));
  OAI21_X1  g216(.A(169), .B1(n287), .B2(n285), .ZN(n288));
  OR3_X1    g217(.A1(n287), .A2(n285), .A3(n194), .ZN(n289));
  AOI21_X1  g218(.A(n282), .B1(n289), .B2(n288), .ZN(n290));
  OR3_X1    g219(.A1(n287), .A2(n285), .A3(n144), .ZN(n291));
  OAI21_X1  g220(.A(200), .B1(n287), .B2(n285), .ZN(n292));
  AND3_X1   g221(.A1(n292), .A2(n291), .A3(n282), .ZN(n293));
  OR2_X1    g222(.A1(n293), .A2(n290), .ZN(n294));
  NAND3_X1  g223(.A1(50), .A2(n120), .A3(n80), .ZN(n295));
  OAI221_X1 g224(.A(n295), .B1(n88), .B2(n157), .C1(68), .C2(n80), .ZN(n296));
  NOR4_X1   g225(.A1(n227), .A2(n147), .A3(n83), .A4(n150), .ZN(n297));
  AOI221_X1 g226(.A(n297), .B1(n150), .B2(n83), .C1(n147), .C2(n296), .ZN(n298));
  NAND3_X1  g227(.A1(349), .A2(232), .A3(n120), .ZN(n299));
  AOI22_X1  g228(.A1(226), .A2(n132), .B1(97), .B2(33), .ZN(n300));
  AOI21_X1  g229(.A(n130), .B1(n300), .B2(n299), .ZN(n301));
  OAI221_X1 g230(.A(238), .B1(n115), .B2(n137), .C1(\1 ), .C2(n235), .ZN(n302));
  OAI21_X1  g231(.A(n302), .B1(n234), .B2(n138), .ZN(n303));
  OAI21_X1  g232(.A(169), .B1(n303), .B2(n301), .ZN(n304));
  NOR3_X1   g233(.A1(n164), .A2(n261), .A3(33), .ZN(n305));
  OAI22_X1  g234(.A1(n84), .A2(n167), .B1(n74), .B2(n120), .ZN(n306));
  OAI21_X1  g235(.A(n163), .B1(n306), .B2(n305), .ZN(n307));
  AOI221_X1 g236(.A(n85), .B1(n128), .B2(n129), .C1(n79), .C2(n233), .ZN(n308));
  AOI21_X1  g237(.A(n308), .B1(n260), .B2(n259), .ZN(n309));
  NAND3_X1  g238(.A1(n309), .A2(n307), .A3(179), .ZN(n310));
  AOI21_X1  g239(.A(n298), .B1(n310), .B2(n304), .ZN(n311));
  NOR3_X1   g240(.A1(n82), .A2(33), .A3(20), .ZN(n312));
  AOI221_X1 g241(.A(n312), .B1(77), .B2(n201), .C1(n83), .C2(20), .ZN(n313));
  NAND4_X1  g242(.A1(n251), .A2(n117), .A3(68), .A4(n124), .ZN(n314));
  OAI221_X1 g243(.A(n314), .B1(n124), .B2(68), .C1(n117), .C2(n313), .ZN(n315));
  NOR3_X1   g244(.A1(n303), .A2(n301), .A3(n144), .ZN(n316));
  AOI21_X1  g245(.A(n146), .B1(n309), .B2(n307), .ZN(n317));
  NOR3_X1   g246(.A1(n317), .A2(n316), .A3(n315), .ZN(n318));
  OR2_X1    g247(.A1(n318), .A2(n311), .ZN(n319));
  OR4_X1    g248(.A1(n294), .A2(n278), .A3(n244), .A4(n319), .ZN(n320));
  NOR2_X1   g249(.A1(n320), .A2(n223), .ZN(4028));
  NAND2_X1  g250(.A1(n214), .A2(n212), .ZN(n322));
  NOR2_X1   g251(.A1(n196), .A2(n193), .ZN(n323));
  NOR4_X1   g252(.A1(n323), .A2(n180), .A3(n155), .A4(n221), .ZN(n324));
  AND2_X1   g253(.A1(n177), .A2(n175), .ZN(n325));
  OAI211_X1 g254(.A(n143), .B(n141), .C1(n155), .C2(n325), .ZN(n326));
  AOI211_X1 g255(.A(n324), .B(n326), .C1(n322), .C2(n181), .ZN(n327));
  INV_X1    g256(.A(n311), .ZN(n328));
  OR3_X1    g257(.A1(n328), .A2(n278), .A3(n244), .ZN(n329));
  AND3_X1   g258(.A1(n290), .A2(n243), .A3(n241), .ZN(n330));
  NOR2_X1   g259(.A1(n319), .A2(n278), .ZN(n331));
  OAI21_X1  g260(.A(n241), .B1(n271), .B2(n244), .ZN(n332));
  AOI21_X1  g261(.A(n332), .B1(n331), .B2(n330), .ZN(n333));
  OAI211_X1 g262(.A(n329), .B(n333), .C1(n327), .C2(n320), .ZN(4145));
  INV_X1    g263(.A(213), .ZN(n335));
  NOR4_X1   g264(.A1(20), .A2(n149), .A3(\1 ), .A4(n335), .ZN(n336));
  NAND2_X1  g265(.A1(n336), .A2(343), .ZN(n337));
  NOR2_X1   g266(.A1(n337), .A2(n219), .ZN(n338));
  XOR2_X1   g267(.A(n338), .B(n221), .ZN(n339));
  INV_X1    g268(.A(n339), .ZN(n340));
  AND2_X1   g269(.A1(n337), .A2(n197), .ZN(n341));
  AOI22_X1  g270(.A1(n340), .A2(n341), .B1(n337), .B2(n322), .ZN(n342));
  INV_X1    g271(.A(330), .ZN(n343));
  NOR2_X1   g272(.A1(n200), .A2(n197), .ZN(n344));
  NOR2_X1   g273(.A1(n337), .A2(n186), .ZN(n345));
  XNOR2_X1  g274(.A(n345), .B(n344), .ZN(n346));
  OR3_X1    g275(.A1(n346), .A2(n339), .A3(n343), .ZN(n347));
  NAND2_X1  g276(.A1(n347), .A2(n342), .ZN(4589));
  INV_X1    g277(.A(n337), .ZN(n349));
  OR2_X1    g278(.A1(n349), .A2(n327), .ZN(n350));
  NOR2_X1   g279(.A1(n174), .A2(179), .ZN(n351));
  NOR3_X1   g280(.A1(n213), .A2(n192), .A3(n142), .ZN(n352));
  NOR4_X1   g281(.A1(n195), .A2(n176), .A3(n140), .A4(n211), .ZN(n353));
  AOI21_X1  g282(.A(n353), .B1(n352), .B2(n351), .ZN(n354));
  MUX2_X1   g283(.S(n337), .B(n223), .A(n354), .ZN(n355));
  OR2_X1    g284(.A1(n355), .A2(n343), .ZN(n356));
  AND2_X1   g285(.A1(n356), .A2(n350), .ZN(n357));
  NOR4_X1   g286(.A1(n80), .A2(13), .A3(n79), .A4(41), .ZN(n358));
  NOR4_X1   g287(.A1(107), .A2(97), .A3(87), .A4(116), .ZN(n359));
  INV_X1    g288(.A(n359), .ZN(n360));
  OR3_X1    g289(.A1(n360), .A2(n358), .A3(n79), .ZN(n361));
  NAND2_X1  g290(.A1(n358), .A2(n96), .ZN(n362));
  OAI211_X1 g291(.A(n361), .B(n362), .C1(n357), .C2(\1 ), .ZN(4667));
  NOR3_X1   g292(.A1(n136), .A2(20), .A3(n149), .ZN(n364));
  NOR2_X1   g293(.A1(n364), .A2(n79), .ZN(n365));
  INV_X1    g294(.A(n365), .ZN(n366));
  XNOR2_X1  g295(.A(n346), .B(330), .ZN(n367));
  NAND2_X1  g296(.A1(n367), .A2(n366), .ZN(n368));
  NOR3_X1   g297(.A1(33), .A2(20), .A3(13), .ZN(n369));
  NAND2_X1  g298(.A1(n369), .A2(n346), .ZN(n370));
  AOI21_X1  g299(.A(n115), .B1(n156), .B2(20), .ZN(n371));
  NOR4_X1   g300(.A1(190), .A2(n194), .A3(n80), .A4(200), .ZN(n372));
  INV_X1    g301(.A(n372), .ZN(n373));
  AND4_X1   g302(.A1(190), .A2(179), .A3(20), .A4(200), .ZN(n374));
  NOR4_X1   g303(.A1(n144), .A2(n194), .A3(n80), .A4(200), .ZN(n375));
  AOI22_X1  g304(.A1(n374), .A2(50), .B1(58), .B2(n375), .ZN(n376));
  OAI21_X1  g305(.A(n376), .B1(n373), .B2(n88), .ZN(n377));
  OAI21_X1  g306(.A(20), .B1(200), .B2(179), .ZN(n378));
  NAND3_X1  g307(.A1(n378), .A2(n144), .A3(20), .ZN(n379));
  OAI21_X1  g308(.A(n120), .B1(n379), .B2(n247), .ZN(n380));
  NAND4_X1  g309(.A1(190), .A2(n194), .A3(20), .A4(200), .ZN(n381));
  OAI21_X1  g310(.A(n378), .B1(190), .B2(n80), .ZN(n382));
  OAI22_X1  g311(.A1(n381), .A2(n73), .B1(n74), .B2(n382), .ZN(n383));
  NOR4_X1   g312(.A1(190), .A2(n194), .A3(n80), .A4(n146), .ZN(n384));
  AND2_X1   g313(.A1(n384), .A2(68), .ZN(n385));
  NAND4_X1  g314(.A1(n144), .A2(n194), .A3(20), .A4(200), .ZN(n386));
  NOR2_X1   g315(.A1(n386), .A2(n75), .ZN(n387));
  OR4_X1    g316(.A1(n385), .A2(n383), .A3(n380), .A4(n387), .ZN(n388));
  INV_X1    g317(.A(311), .ZN(n389));
  AOI22_X1  g318(.A1(n374), .A2(326), .B1(322), .B2(n375), .ZN(n390));
  OAI21_X1  g319(.A(n390), .B1(n373), .B2(n389), .ZN(n391));
  NAND4_X1  g320(.A1(329), .A2(n144), .A3(20), .A4(n378), .ZN(n392));
  NAND2_X1  g321(.A1(n392), .A2(33), .ZN(n393));
  OAI22_X1  g322(.A1(n381), .A2(n188), .B1(n207), .B2(n382), .ZN(n394));
  INV_X1    g323(.A(317), .ZN(n395));
  INV_X1    g324(.A(n384), .ZN(n396));
  OAI22_X1  g325(.A1(n396), .A2(n395), .B1(n166), .B2(n386), .ZN(n397));
  OR4_X1    g326(.A1(n394), .A2(n393), .A3(n391), .A4(n397), .ZN(n398));
  OAI21_X1  g327(.A(n398), .B1(n388), .B2(n377), .ZN(n399));
  NOR4_X1   g328(.A1(n80), .A2(13), .A3(n79), .A4(n120), .ZN(n400));
  OAI211_X1 g329(.A(50), .B(n136), .C1(58), .C2(68), .ZN(n401));
  OAI211_X1 g330(.A(n400), .B(n401), .C1(n113), .C2(n136), .ZN(n402));
  NOR4_X1   g331(.A1(n80), .A2(13), .A3(n79), .A4(33), .ZN(n403));
  NAND3_X1  g332(.A1(20), .A2(n149), .A3(\1 ), .ZN(n404));
  AOI22_X1  g333(.A1(n403), .A2(1947), .B1(n182), .B2(n404), .ZN(n405));
  NOR2_X1   g334(.A1(n371), .A2(n369), .ZN(n406));
  INV_X1    g335(.A(n406), .ZN(n407));
  AOI21_X1  g336(.A(n407), .B1(n405), .B2(n402), .ZN(n408));
  NOR3_X1   g337(.A1(n364), .A2(n358), .A3(n79), .ZN(n409));
  INV_X1    g338(.A(n409), .ZN(n410));
  AOI211_X1 g339(.A(n408), .B(n410), .C1(n399), .C2(n371), .ZN(n411));
  AOI22_X1  g340(.A1(n370), .A2(n411), .B1(n367), .B2(n358), .ZN(n412));
  NAND2_X1  g341(.A1(n412), .A2(n368), .ZN(4815));
  NOR2_X1   g342(.A1(n337), .A2(n282), .ZN(n414));
  XOR2_X1   g343(.A(n414), .B(n294), .ZN(n415));
  XNOR2_X1  g344(.A(n415), .B(n350), .ZN(n416));
  XNOR2_X1  g345(.A(n416), .B(n356), .ZN(n417));
  XOR2_X1   g346(.A(n416), .B(n356), .ZN(n418));
  NOR2_X1   g347(.A1(33), .A2(13), .ZN(n419));
  NAND2_X1  g348(.A1(n419), .A2(n415), .ZN(n420));
  INV_X1    g349(.A(n371), .ZN(n421));
  AOI22_X1  g350(.A1(n374), .A2(137), .B1(143), .B2(n375), .ZN(n422));
  OAI21_X1  g351(.A(n422), .B1(n373), .B2(n247), .ZN(n423));
  INV_X1    g352(.A(132), .ZN(n424));
  OAI21_X1  g353(.A(n120), .B1(n379), .B2(n424), .ZN(n425));
  OAI22_X1  g354(.A1(n381), .A2(n82), .B1(n95), .B2(n382), .ZN(n426));
  INV_X1    g355(.A(150), .ZN(n427));
  OAI22_X1  g356(.A1(n396), .A2(n427), .B1(n83), .B2(n386), .ZN(n428));
  OR4_X1    g357(.A1(n426), .A2(n425), .A3(n423), .A4(n428), .ZN(n429));
  AOI22_X1  g358(.A1(n374), .A2(303), .B1(294), .B2(n375), .ZN(n430));
  OAI21_X1  g359(.A(n430), .B1(n373), .B2(n182), .ZN(n431));
  OAI21_X1  g360(.A(33), .B1(n379), .B2(n389), .ZN(n432));
  OAI22_X1  g361(.A1(n381), .A2(n75), .B1(n74), .B2(n382), .ZN(n433));
  OAI22_X1  g362(.A1(n396), .A2(n166), .B1(n73), .B2(n386), .ZN(n434));
  OR4_X1    g363(.A1(n433), .A2(n432), .A3(n431), .A4(n434), .ZN(n435));
  AOI21_X1  g364(.A(n421), .B1(n435), .B2(n429), .ZN(n436));
  NOR2_X1   g365(.A1(n419), .A2(n371), .ZN(n437));
  AOI211_X1 g366(.A(n436), .B(n410), .C1(n88), .C2(n437), .ZN(n438));
  AOI22_X1  g367(.A1(n420), .A2(n438), .B1(n418), .B2(n358), .ZN(n439));
  OAI21_X1  g368(.A(n439), .B1(n417), .B2(n365), .ZN(4944));
  NAND2_X1  g369(.A1(n149), .A2(\1 ), .ZN(n441));
  NOR2_X1   g370(.A1(n318), .A2(n311), .ZN(n442));
  NOR2_X1   g371(.A1(n337), .A2(n298), .ZN(n443));
  XNOR2_X1  g372(.A(n443), .B(n442), .ZN(n444));
  INV_X1    g373(.A(n336), .ZN(n445));
  NOR2_X1   g374(.A1(n445), .A2(n274), .ZN(n446));
  XOR2_X1   g375(.A(n446), .B(n278), .ZN(n447));
  OR4_X1    g376(.A1(n444), .A2(n415), .A3(n355), .A4(n447), .ZN(n448));
  NOR2_X1   g377(.A1(n355), .A2(n320), .ZN(n449));
  XNOR2_X1  g378(.A(n449), .B(n448), .ZN(n450));
  NAND2_X1  g379(.A1(n450), .A2(330), .ZN(n451));
  OR3_X1    g380(.A1(n349), .A2(n327), .A3(n320), .ZN(n452));
  NAND3_X1  g381(.A1(n452), .A2(n333), .A3(n329), .ZN(n453));
  OR2_X1    g382(.A1(n447), .A2(n444), .ZN(n454));
  NOR4_X1   g383(.A1(n415), .A2(n349), .A3(n327), .A4(n454), .ZN(n455));
  AOI211_X1 g384(.A(n282), .B(n349), .C1(n289), .C2(n288), .ZN(n456));
  INV_X1    g385(.A(n456), .ZN(n457));
  OAI211_X1 g386(.A(n253), .B(n445), .C1(n270), .C2(n264), .ZN(n458));
  AOI211_X1 g387(.A(n298), .B(n349), .C1(n310), .C2(n304), .ZN(n459));
  INV_X1    g388(.A(n459), .ZN(n460));
  OAI221_X1 g389(.A(n458), .B1(n457), .B2(n454), .C1(n447), .C2(n460), .ZN(n461));
  NOR2_X1   g390(.A1(n461), .A2(n455), .ZN(n462));
  XOR2_X1   g391(.A(n462), .B(n453), .ZN(n463));
  XNOR2_X1  g392(.A(n463), .B(n451), .ZN(n464));
  AOI21_X1  g393(.A(n79), .B1(n80), .B2(13), .ZN(n465));
  AND2_X1   g394(.A1(77), .A2(50), .ZN(n466));
  AOI22_X1  g395(.A1(n245), .A2(n466), .B1(68), .B2(n82), .ZN(n467));
  NAND3_X1  g396(.A1(n158), .A2(n78), .A3(116), .ZN(n468));
  OAI221_X1 g397(.A(n468), .B1(n465), .B2(n464), .C1(n441), .C2(n467), .ZN(5002));
  INV_X1    g398(.A(n358), .ZN(n470));
  NOR2_X1   g399(.A1(n337), .A2(n162), .ZN(n471));
  XOR2_X1   g400(.A(n471), .B(n180), .ZN(n472));
  OR4_X1    g401(.A1(n346), .A2(n339), .A3(n343), .A4(n472), .ZN(n473));
  NOR2_X1   g402(.A1(n337), .A2(n153), .ZN(n474));
  XOR2_X1   g403(.A(n474), .B(n155), .ZN(n475));
  NOR4_X1   g404(.A1(n339), .A2(n349), .A3(n323), .A4(n472), .ZN(n476));
  NAND2_X1  g405(.A1(n337), .A2(n322), .ZN(n477));
  OAI22_X1  g406(.A1(n477), .A2(n472), .B1(n349), .B2(n325), .ZN(n478));
  NOR2_X1   g407(.A1(n478), .A2(n476), .ZN(n479));
  XNOR2_X1  g408(.A(n479), .B(n475), .ZN(n480));
  XNOR2_X1  g409(.A(n480), .B(n473), .ZN(n481));
  XNOR2_X1  g410(.A(n472), .B(n342), .ZN(n482));
  XOR2_X1   g411(.A(n482), .B(n347), .ZN(n483));
  OR2_X1    g412(.A1(n346), .A2(n343), .ZN(n484));
  XOR2_X1   g413(.A(n341), .B(n339), .ZN(n485));
  XNOR2_X1  g414(.A(n485), .B(n484), .ZN(n486));
  INV_X1    g415(.A(n486), .ZN(n487));
  NAND3_X1  g416(.A1(n487), .A2(n483), .A3(n357), .ZN(n488));
  AOI211_X1 g417(.A(n481), .B(n470), .C1(n357), .C2(n488), .ZN(n489));
  NAND2_X1  g418(.A1(n475), .A2(n369), .ZN(n490));
  AOI22_X1  g419(.A1(n374), .A2(143), .B1(150), .B2(n375), .ZN(n491));
  OAI21_X1  g420(.A(n491), .B1(n373), .B2(n82), .ZN(n492));
  INV_X1    g421(.A(137), .ZN(n493));
  OAI21_X1  g422(.A(n120), .B1(n379), .B2(n493), .ZN(n494));
  OAI22_X1  g423(.A1(n381), .A2(n95), .B1(n83), .B2(n382), .ZN(n495));
  OAI22_X1  g424(.A1(n396), .A2(n247), .B1(n88), .B2(n386), .ZN(n496));
  OR4_X1    g425(.A1(n495), .A2(n494), .A3(n492), .A4(n496), .ZN(n497));
  AOI22_X1  g426(.A1(n374), .A2(311), .B1(303), .B2(n375), .ZN(n498));
  OAI21_X1  g427(.A(n498), .B1(n373), .B2(n166), .ZN(n499));
  OAI21_X1  g428(.A(33), .B1(n379), .B2(n395), .ZN(n500));
  OAI22_X1  g429(.A1(n381), .A2(n182), .B1(n75), .B2(n382), .ZN(n501));
  OAI22_X1  g430(.A1(n396), .A2(n207), .B1(n74), .B2(n386), .ZN(n502));
  OR4_X1    g431(.A1(n501), .A2(n500), .A3(n499), .A4(n502), .ZN(n503));
  AOI21_X1  g432(.A(n421), .B1(n503), .B2(n497), .ZN(n504));
  INV_X1    g433(.A(n400), .ZN(n505));
  AOI21_X1  g434(.A(n403), .B1(n404), .B2(n73), .ZN(n506));
  OAI21_X1  g435(.A(n506), .B1(n505), .B2(n103), .ZN(n507));
  AOI211_X1 g436(.A(n504), .B(n410), .C1(n406), .C2(n507), .ZN(n508));
  NAND2_X1  g437(.A1(n508), .A2(n490), .ZN(n509));
  OAI21_X1  g438(.A(n509), .B1(n481), .B2(n365), .ZN(n510));
  NOR2_X1   g439(.A1(n510), .A2(n489), .ZN(n511));
  INV_X1    g440(.A(n511), .ZN(5045));
  AND2_X1   g441(.A1(n487), .A2(n357), .ZN(n513));
  OAI21_X1  g442(.A(n358), .B1(n487), .B2(n357), .ZN(n514));
  AND2_X1   g443(.A1(n369), .A2(n339), .ZN(n515));
  AND2_X1   g444(.A1(n374), .A2(159), .ZN(n516));
  AOI221_X1 g445(.A(n516), .B1(n372), .B2(68), .C1(50), .C2(n375), .ZN(n517));
  OAI21_X1  g446(.A(n120), .B1(n386), .B2(n74), .ZN(n518));
  OAI22_X1  g447(.A1(n381), .A2(n88), .B1(n73), .B2(n382), .ZN(n519));
  OAI22_X1  g448(.A1(n379), .A2(n427), .B1(n95), .B2(n396), .ZN(n520));
  NOR3_X1   g449(.A1(n520), .A2(n519), .A3(n518), .ZN(n521));
  AOI22_X1  g450(.A1(n374), .A2(322), .B1(317), .B2(n375), .ZN(n522));
  OAI21_X1  g451(.A(n522), .B1(n373), .B2(n188), .ZN(n523));
  NAND4_X1  g452(.A1(326), .A2(n144), .A3(20), .A4(n378), .ZN(n524));
  NAND2_X1  g453(.A1(n524), .A2(33), .ZN(n525));
  OAI22_X1  g454(.A1(n381), .A2(n207), .B1(n166), .B2(n382), .ZN(n526));
  OAI22_X1  g455(.A1(n396), .A2(n389), .B1(n182), .B2(n386), .ZN(n527));
  NOR4_X1   g456(.A1(n526), .A2(n525), .A3(n523), .A4(n527), .ZN(n528));
  AOI21_X1  g457(.A(n528), .B1(n521), .B2(n517), .ZN(n529));
  AND2_X1   g458(.A1(77), .A2(68), .ZN(n530));
  NOR4_X1   g459(.A1(n95), .A2(50), .A3(45), .A4(n530), .ZN(n531));
  AOI221_X1 g460(.A(n505), .B1(n359), .B2(n531), .C1(n106), .C2(45), .ZN(n532));
  AOI221_X1 g461(.A(n532), .B1(n403), .B2(n360), .C1(n75), .C2(n404), .ZN(n533));
  OAI221_X1 g462(.A(n409), .B1(n407), .B2(n533), .C1(n421), .C2(n529), .ZN(n534));
  OR2_X1    g463(.A1(n534), .A2(n515), .ZN(n535));
  OAI221_X1 g464(.A(n535), .B1(n513), .B2(n514), .C1(n486), .C2(n365), .ZN(5047));
  XNOR2_X1  g465(.A(n513), .B(n483), .ZN(n537));
  NAND2_X1  g466(.A1(n472), .A2(n369), .ZN(n538));
  AOI22_X1  g467(.A1(n374), .A2(150), .B1(159), .B2(n375), .ZN(n539));
  OAI21_X1  g468(.A(n539), .B1(n373), .B2(n95), .ZN(n540));
  OAI21_X1  g469(.A(n120), .B1(n386), .B2(n73), .ZN(n541));
  OAI22_X1  g470(.A1(n381), .A2(n83), .B1(n88), .B2(n382), .ZN(n542));
  INV_X1    g471(.A(143), .ZN(n543));
  OAI22_X1  g472(.A1(n379), .A2(n543), .B1(n82), .B2(n396), .ZN(n544));
  OR4_X1    g473(.A1(n542), .A2(n541), .A3(n540), .A4(n544), .ZN(n545));
  AOI22_X1  g474(.A1(n374), .A2(317), .B1(311), .B2(n375), .ZN(n546));
  OAI21_X1  g475(.A(n546), .B1(n373), .B2(n207), .ZN(n547));
  OAI22_X1  g476(.A1(n381), .A2(n166), .B1(n182), .B2(n382), .ZN(n548));
  NAND4_X1  g477(.A1(322), .A2(n144), .A3(20), .A4(n378), .ZN(n549));
  OAI21_X1  g478(.A(n549), .B1(n396), .B2(n188), .ZN(n550));
  OR4_X1    g479(.A1(n548), .A2(n387), .A3(n120), .A4(n550), .ZN(n551));
  OAI21_X1  g480(.A(n545), .B1(n551), .B2(n547), .ZN(n552));
  AOI21_X1  g481(.A(n403), .B1(n404), .B2(n74), .ZN(n553));
  OAI21_X1  g482(.A(n553), .B1(n505), .B2(n110), .ZN(n554));
  AOI221_X1 g483(.A(n410), .B1(n406), .B2(n554), .C1(n371), .C2(n552), .ZN(n555));
  AOI22_X1  g484(.A1(n538), .A2(n555), .B1(n483), .B2(n366), .ZN(n556));
  OAI21_X1  g485(.A(n556), .B1(n537), .B2(n470), .ZN(5078));
  NOR4_X1   g486(.A1(n415), .A2(n355), .A3(n343), .A4(n444), .ZN(n558));
  INV_X1    g487(.A(n447), .ZN(n559));
  OR4_X1    g488(.A1(n415), .A2(n349), .A3(n327), .A4(n444), .ZN(n560));
  XOR2_X1   g489(.A(n443), .B(n442), .ZN(n561));
  AOI21_X1  g490(.A(n459), .B1(n456), .B2(n561), .ZN(n562));
  NAND3_X1  g491(.A1(n562), .A2(n560), .A3(n559), .ZN(n563));
  NOR4_X1   g492(.A1(n415), .A2(n349), .A3(n327), .A4(n444), .ZN(n564));
  OAI21_X1  g493(.A(n460), .B1(n457), .B2(n444), .ZN(n565));
  OAI21_X1  g494(.A(n447), .B1(n565), .B2(n564), .ZN(n566));
  AND2_X1   g495(.A1(n566), .A2(n563), .ZN(n567));
  XNOR2_X1  g496(.A(n567), .B(n558), .ZN(n568));
  OR3_X1    g497(.A1(n415), .A2(n355), .A3(n343), .ZN(n569));
  NOR3_X1   g498(.A1(n415), .A2(n349), .A3(n327), .ZN(n570));
  NOR3_X1   g499(.A1(n570), .A2(n456), .A3(n444), .ZN(n571));
  OR3_X1    g500(.A1(n415), .A2(n349), .A3(n327), .ZN(n572));
  AOI21_X1  g501(.A(n561), .B1(n572), .B2(n457), .ZN(n573));
  OR3_X1    g502(.A1(n573), .A2(n571), .A3(n569), .ZN(n574));
  OAI21_X1  g503(.A(n569), .B1(n573), .B2(n571), .ZN(n575));
  OR3_X1    g504(.A1(n355), .A2(n320), .A3(n343), .ZN(n576));
  NAND4_X1  g505(.A1(n452), .A2(n333), .A3(n329), .A4(n576), .ZN(n577));
  AOI21_X1  g506(.A(n577), .B1(n575), .B2(n574), .ZN(n578));
  XNOR2_X1  g507(.A(n578), .B(n568), .ZN(n579));
  INV_X1    g508(.A(n437), .ZN(n580));
  AOI22_X1  g509(.A1(n374), .A2(128), .B1(132), .B2(n375), .ZN(n581));
  OAI21_X1  g510(.A(n581), .B1(n373), .B2(n543), .ZN(n582));
  NAND4_X1  g511(.A1(n144), .A2(125), .A3(20), .A4(n378), .ZN(n583));
  NAND2_X1  g512(.A1(n583), .A2(n120), .ZN(n584));
  OAI22_X1  g513(.A1(n381), .A2(n427), .B1(n247), .B2(n382), .ZN(n585));
  OAI22_X1  g514(.A1(n396), .A2(n493), .B1(n82), .B2(n386), .ZN(n586));
  NOR4_X1   g515(.A1(n585), .A2(n584), .A3(n582), .A4(n586), .ZN(n587));
  AND2_X1   g516(.A1(n374), .A2(283), .ZN(n588));
  AOI221_X1 g517(.A(n588), .B1(n372), .B2(97), .C1(116), .C2(n375), .ZN(n589));
  OAI21_X1  g518(.A(33), .B1(n386), .B2(n83), .ZN(n590));
  OAI22_X1  g519(.A1(n381), .A2(n73), .B1(n88), .B2(n382), .ZN(n591));
  OAI22_X1  g520(.A1(n379), .A2(n207), .B1(n75), .B2(n396), .ZN(n592));
  NOR3_X1   g521(.A1(n592), .A2(n591), .A3(n590), .ZN(n593));
  AOI21_X1  g522(.A(n587), .B1(n593), .B2(n589), .ZN(n594));
  OAI221_X1 g523(.A(n409), .B1(n421), .B2(n594), .C1(58), .C2(n580), .ZN(n595));
  AOI21_X1  g524(.A(n595), .B1(n447), .B2(n419), .ZN(n596));
  AOI21_X1  g525(.A(n596), .B1(n568), .B2(n366), .ZN(n597));
  OAI21_X1  g526(.A(n597), .B1(n579), .B2(n470), .ZN(5102));
  NOR2_X1   g527(.A1(n445), .A2(n229), .ZN(n599));
  XOR2_X1   g528(.A(n599), .B(n244), .ZN(n600));
  NOR3_X1   g529(.A1(n600), .A2(n461), .A3(n455), .ZN(n601));
  OR4_X1    g530(.A1(n415), .A2(n349), .A3(n327), .A4(n454), .ZN(n602));
  NOR3_X1   g531(.A1(n457), .A2(n447), .A3(n444), .ZN(n603));
  OAI21_X1  g532(.A(n458), .B1(n460), .B2(n447), .ZN(n604));
  NOR2_X1   g533(.A1(n604), .A2(n603), .ZN(n605));
  XNOR2_X1  g534(.A(n599), .B(n244), .ZN(n606));
  AOI21_X1  g535(.A(n606), .B1(n605), .B2(n602), .ZN(n607));
  NOR4_X1   g536(.A1(n601), .A2(n448), .A3(n343), .A4(n607), .ZN(n608));
  NOR4_X1   g537(.A1(n444), .A2(n415), .A3(n355), .A4(n447), .ZN(n609));
  NAND3_X1  g538(.A1(n606), .A2(n605), .A3(n602), .ZN(n610));
  OAI21_X1  g539(.A(n600), .B1(n461), .B2(n455), .ZN(n611));
  AOI22_X1  g540(.A1(n610), .A2(n611), .B1(n609), .B2(330), .ZN(n612));
  OR2_X1    g541(.A1(n612), .A2(n608), .ZN(n613));
  NOR3_X1   g542(.A1(n573), .A2(n571), .A3(n569), .ZN(n614));
  NOR3_X1   g543(.A1(n415), .A2(n355), .A3(n343), .ZN(n615));
  NAND3_X1  g544(.A1(n572), .A2(n457), .A3(n561), .ZN(n616));
  OAI21_X1  g545(.A(n444), .B1(n570), .B2(n456), .ZN(n617));
  AOI21_X1  g546(.A(n615), .B1(n617), .B2(n616), .ZN(n618));
  AOI21_X1  g547(.A(n453), .B1(n449), .B2(330), .ZN(n619));
  OAI21_X1  g548(.A(n619), .B1(n618), .B2(n614), .ZN(n620));
  OAI21_X1  g549(.A(n577), .B1(n612), .B2(n608), .ZN(n621));
  AND3_X1   g550(.A1(n566), .A2(n563), .A3(n558), .ZN(n622));
  AOI21_X1  g551(.A(n558), .B1(n566), .B2(n563), .ZN(n623));
  OAI22_X1  g552(.A1(n608), .A2(n612), .B1(n623), .B2(n622), .ZN(n624));
  OAI21_X1  g553(.A(n621), .B1(n624), .B2(n620), .ZN(n625));
  NOR2_X1   g554(.A1(41), .A2(33), .ZN(n626));
  INV_X1    g555(.A(n626), .ZN(n627));
  NAND2_X1  g556(.A1(n374), .A2(125), .ZN(n628));
  AOI22_X1  g557(.A1(n375), .A2(128), .B1(132), .B2(n384), .ZN(n629));
  NAND2_X1  g558(.A1(n629), .A2(n628), .ZN(n630));
  OAI21_X1  g559(.A(n626), .B1(n386), .B2(n247), .ZN(n631));
  NAND4_X1  g560(.A1(n144), .A2(124), .A3(20), .A4(n378), .ZN(n632));
  OAI21_X1  g561(.A(n632), .B1(n382), .B2(n427), .ZN(n633));
  OAI22_X1  g562(.A1(n373), .A2(n493), .B1(n543), .B2(n381), .ZN(n634));
  NOR4_X1   g563(.A1(n633), .A2(n631), .A3(n630), .A4(n634), .ZN(n635));
  AOI21_X1  g564(.A(50), .B1(n170), .B2(33), .ZN(n636));
  AND2_X1   g565(.A1(n374), .A2(116), .ZN(n637));
  AOI221_X1 g566(.A(n637), .B1(n375), .B2(107), .C1(97), .C2(n384), .ZN(n638));
  OAI211_X1 g567(.A(n170), .B(33), .C1(n95), .C2(n386), .ZN(n639));
  OAI22_X1  g568(.A1(n379), .A2(n166), .B1(n83), .B2(n382), .ZN(n640));
  OAI22_X1  g569(.A1(n373), .A2(n73), .B1(n88), .B2(n381), .ZN(n641));
  NOR3_X1   g570(.A1(n641), .A2(n640), .A3(n639), .ZN(n642));
  AOI221_X1 g571(.A(n635), .B1(n636), .B2(n627), .C1(n642), .C2(n638), .ZN(n643));
  OAI221_X1 g572(.A(n409), .B1(n421), .B2(n643), .C1(50), .C2(n580), .ZN(n644));
  AOI21_X1  g573(.A(n644), .B1(n600), .B2(n419), .ZN(n645));
  AOI221_X1 g574(.A(n645), .B1(n613), .B2(n366), .C1(n358), .C2(n625), .ZN(n646));
  INV_X1    g575(.A(n646), .ZN(5120));
  NOR3_X1   g576(.A1(n619), .A2(n618), .A3(n614), .ZN(n648));
  OR3_X1    g577(.A1(n648), .A2(n578), .A3(n470), .ZN(n649));
  NOR2_X1   g578(.A1(n573), .A2(n571), .ZN(n650));
  XNOR2_X1  g579(.A(n650), .B(n615), .ZN(n651));
  AND2_X1   g580(.A1(n374), .A2(132), .ZN(n652));
  AOI221_X1 g581(.A(n652), .B1(n372), .B2(150), .C1(137), .C2(n375), .ZN(n653));
  OAI21_X1  g582(.A(n120), .B1(n386), .B2(n95), .ZN(n654));
  OAI22_X1  g583(.A1(n381), .A2(n247), .B1(n82), .B2(n382), .ZN(n655));
  AND2_X1   g584(.A1(n384), .A2(143), .ZN(n656));
  AND4_X1   g585(.A1(n144), .A2(128), .A3(20), .A4(n378), .ZN(n657));
  NOR4_X1   g586(.A1(n656), .A2(n655), .A3(n654), .A4(n657), .ZN(n658));
  AND2_X1   g587(.A1(n374), .A2(294), .ZN(n659));
  AOI221_X1 g588(.A(n659), .B1(n372), .B2(107), .C1(283), .C2(n375), .ZN(n660));
  OAI21_X1  g589(.A(33), .B1(n386), .B2(n88), .ZN(n661));
  OAI22_X1  g590(.A1(n381), .A2(n74), .B1(n73), .B2(n382), .ZN(n662));
  OAI22_X1  g591(.A1(n379), .A2(n188), .B1(n182), .B2(n396), .ZN(n663));
  NOR3_X1   g592(.A1(n663), .A2(n662), .A3(n661), .ZN(n664));
  AOI22_X1  g593(.A1(n660), .A2(n664), .B1(n658), .B2(n653), .ZN(n665));
  OAI221_X1 g594(.A(n409), .B1(n421), .B2(n665), .C1(68), .C2(n580), .ZN(n666));
  AOI21_X1  g595(.A(n666), .B1(n444), .B2(n419), .ZN(n667));
  AOI21_X1  g596(.A(n667), .B1(n651), .B2(n366), .ZN(n668));
  AND2_X1   g597(.A1(n668), .A2(n649), .ZN(n669));
  INV_X1    g598(.A(n669), .ZN(5121));
  NOR4_X1   g599(.A1(5047), .A2(4944), .A3(4815), .A4(5078), .ZN(n671));
  NAND4_X1  g600(.A1(n669), .A2(n646), .A3(n511), .A4(n671), .ZN(n672));
  OR2_X1    g601(.A1(n672), .A2(5102), .ZN(5192));
  NOR2_X1   g602(.A1(343), .A2(n335), .ZN(n674));
  NAND2_X1  g603(.A1(n674), .A2(n646), .ZN(n675));
  OAI211_X1 g604(.A(5192), .B(213), .C1(5102), .C2(n675), .ZN(5231));
  XOR2_X1   g605(.A(5078), .B(n511), .ZN(n677));
  XNOR2_X1  g606(.A(5047), .B(4815), .ZN(n678));
  XNOR2_X1  g607(.A(n678), .B(n677), .ZN(n679));
  OAI211_X1 g608(.A(5102), .B(n646), .C1(343), .C2(n335), .ZN(n680));
  OR3_X1    g609(.A1(n674), .A2(n646), .A3(5102), .ZN(n681));
  INV_X1    g610(.A(350), .ZN(n682));
  NOR3_X1   g611(.A1(n682), .A2(343), .A3(n335), .ZN(n683));
  XOR2_X1   g612(.A(n669), .B(4944), .ZN(n684));
  AND4_X1   g613(.A1(n683), .A2(n681), .A3(n680), .A4(n684), .ZN(n685));
  INV_X1    g614(.A(n683), .ZN(n686));
  XNOR2_X1  g615(.A(n669), .B(4944), .ZN(n687));
  AND4_X1   g616(.A1(n686), .A2(n681), .A3(n680), .A4(n687), .ZN(n688));
  AOI211_X1 g617(.A(n683), .B(n687), .C1(n681), .C2(n680), .ZN(n689));
  AOI211_X1 g618(.A(n686), .B(n684), .C1(n681), .C2(n680), .ZN(n690));
  NOR4_X1   g619(.A1(n689), .A2(n688), .A3(n685), .A4(n690), .ZN(n691));
  XNOR2_X1  g620(.A(n691), .B(n679), .ZN(5360));
  XOR2_X1   g621(.A(n646), .B(5102), .ZN(n693));
  XNOR2_X1  g622(.A(n693), .B(n684), .ZN(n694));
  XNOR2_X1  g623(.A(n694), .B(n679), .ZN(5361));
endmodule


