// Benchmark "c2670" written by ABC on Tue Dec 06 12:35:51 2022

module c2670 ( 
    \1 , 2, 3, 4, 5, 6, 7, 8, 11, 14, 15, 16, 19, 20, 21, 22, 23, 24, 25,
    26, 27, 28, 29, 32, 33, 34, 35, 36, 37, 40, 43, 44, 47, 48, 49, 50, 51,
    52, 53, 54, 55, 56, 57, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 72, 73,
    74, 75, 76, 77, 78, 79, 80, 81, 82, 85, 86, 87, 88, 89, 90, 91, 92, 93,
    94, 95, 96, 99, 100, 101, 102, 103, 104, 105, 106, 107, 108, 111, 112,
    113, 114, 115, 116, 117, 118, 119, 120, 123, 124, 125, 126, 127, 128,
    129, 130, 131, 132, 135, 136, 137, 138, 139, 140, 141, 142, 143, 144,
    145, 146, 147, 148, 149, 150, 151, 152, 153, 154, 155, 156, 157, 158,
    159, 160, 161, 162, 163, 164, 165, 166, 167, 168, 169, 170, 171, 172,
    173, 174, 175, 176, 177, 178, 179, 180, 181, 182, 183, 184, 185, 186,
    187, 188, 189, 190, 191, 192, 193, 194, 195, 196, 197, 198, 199, 200,
    201, 202, 203, 204, 205, 206, 207, 208, 209, 210, 211, 212, 213, 214,
    215, 216, 217, 218, 219, 224, 227, 230, 231, 234, 237, 241, 246, 253,
    256, 259, 262, 263, 266, 269, 272, 275, 278, 281, 284, 287, 290, 294,
    297, 301, 305, 309, 313, 316, 319, 322, 325, 328, 331, 334, 337, 340,
    343, 346, 349, 352, 355,
    398, 400, 401, 419, 420, 456, 457, 458, 487, 488, 489, 490, 491, 492,
    493, 494, 792, 799, 805, 1026, 1028, 1029, 1269, 1277, 1448, 1726,
    1816, 1817, 1818, 1819, 1820, 1821, 1969, 1970, 1971, 2010, 2012, 2014,
    2016, 2018, 2020, 2022, 2387, 2388, 2389, 2390, 2496, 2643, 2644, 2891,
    2925, 2970, 2971, 3038, 3079, 3546, 3671, 3803, 3804, 3809, 3851, 3875,
    3881, 3882  );
  input  \1 , 2, 3, 4, 5, 6, 7, 8, 11, 14, 15, 16, 19, 20, 21, 22, 23,
    24, 25, 26, 27, 28, 29, 32, 33, 34, 35, 36, 37, 40, 43, 44, 47, 48, 49,
    50, 51, 52, 53, 54, 55, 56, 57, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69,
    72, 73, 74, 75, 76, 77, 78, 79, 80, 81, 82, 85, 86, 87, 88, 89, 90, 91,
    92, 93, 94, 95, 96, 99, 100, 101, 102, 103, 104, 105, 106, 107, 108,
    111, 112, 113, 114, 115, 116, 117, 118, 119, 120, 123, 124, 125, 126,
    127, 128, 129, 130, 131, 132, 135, 136, 137, 138, 139, 140, 141, 142,
    143, 144, 145, 146, 147, 148, 149, 150, 151, 152, 153, 154, 155, 156,
    157, 158, 159, 160, 161, 162, 163, 164, 165, 166, 167, 168, 169, 170,
    171, 172, 173, 174, 175, 176, 177, 178, 179, 180, 181, 182, 183, 184,
    185, 186, 187, 188, 189, 190, 191, 192, 193, 194, 195, 196, 197, 198,
    199, 200, 201, 202, 203, 204, 205, 206, 207, 208, 209, 210, 211, 212,
    213, 214, 215, 216, 217, 218, 219, 224, 227, 230, 231, 234, 237, 241,
    246, 253, 256, 259, 262, 263, 266, 269, 272, 275, 278, 281, 284, 287,
    290, 294, 297, 301, 305, 309, 313, 316, 319, 322, 325, 328, 331, 334,
    337, 340, 343, 346, 349, 352, 355;
  output 398, 400, 401, 419, 420, 456, 457, 458, 487, 488, 489, 490, 491, 492,
    493, 494, 792, 799, 805, 1026, 1028, 1029, 1269, 1277, 1448, 1726,
    1816, 1817, 1818, 1819, 1820, 1821, 1969, 1970, 1971, 2010, 2012, 2014,
    2016, 2018, 2020, 2022, 2387, 2388, 2389, 2390, 2496, 2643, 2644, 2891,
    2925, 2970, 2971, 3038, 3079, 3546, 3671, 3803, 3804, 3809, 3851, 3875,
    3881, 3882;
  wire n387, n388, n391, n392, n393, n394, n396, n397, n398, n399, n400,
    n401, n402, n404, n405, n406, n407, n409, n410, n411, n412, n414, n415,
    n416, n417, n418, n419, n421, n422, n423, n424, n427, n428, n429, n431,
    n432, n433, n435, n437, n439, n440, n441, n445, n446, n447, n449, n450,
    n451, n452, n454, n455, n456, n457, n459, n460, n461, n462, n463, n464,
    n467, n469, n470, n471, n472, n474, n475, n476, n477, n478, n479, n480,
    n481, n482, n483, n485, n486, n487, n488, n489, n490, n491, n492, n493,
    n494, n495, n496, n497, n498, n499, n501, n502, n503, n504, n505, n506,
    n507, n508, n509, n510, n511, n512, n514, n515, n516, n517, n518, n519,
    n520, n521, n522, n523, n524, n525, n526, n527, n529, n530, n531, n532,
    n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
    n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
    n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
    n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
    n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
    n593, n594, n595, n596, n597, n600, n601, n602, n603, n604, n605, n606,
    n607, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
    n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n631, n632,
    n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n645,
    n646, n647, n648, n649, n650, n651, n652, n654, n655, n656, n657, n658,
    n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
    n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
    n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
    n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
    n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
    n719, n722, n723;
  INV_X1    g000(.A(44), .ZN(487));
  INV_X1    g001(.A(132), .ZN(488));
  INV_X1    g002(.A(82), .ZN(489));
  INV_X1    g003(.A(96), .ZN(490));
  INV_X1    g004(.A(69), .ZN(491));
  INV_X1    g005(.A(120), .ZN(492));
  INV_X1    g006(.A(57), .ZN(493));
  INV_X1    g007(.A(108), .ZN(494));
  NAND4_X1  g008(.A1(305), .A2(301), .A3(297), .A4(309), .ZN(792));
  NAND3_X1  g009(.A1(237), .A2(15), .A3(2), .ZN(799));
  AND2_X1   g010(.A1(219), .A2(94), .ZN(1026));
  NAND2_X1  g011(.A1(237), .A2(7), .ZN(1028));
  NAND3_X1  g012(.A1(237), .A2(231), .A3(7), .ZN(1029));
  NAND3_X1  g013(.A1(325), .A2(237), .A3(7), .ZN(1269));
  AND4_X1   g014(.A1(108), .A2(69), .A3(57), .A4(120), .ZN(n387));
  AND4_X1   g015(.A1(96), .A2(82), .A3(44), .A4(132), .ZN(n388));
  AND2_X1   g016(.A1(n388), .A2(n387), .ZN(1277));
  INV_X1    g017(.A(1277), .ZN(1448));
  INV_X1    g018(.A(325), .ZN(n391));
  NOR2_X1   g019(.A1(n388), .A2(n391), .ZN(n392));
  INV_X1    g020(.A(231), .ZN(n393));
  NOR2_X1   g021(.A1(n387), .A2(n393), .ZN(n394));
  NOR2_X1   g022(.A1(n394), .A2(n392), .ZN(1726));
  NAND3_X1  g023(.A1(322), .A2(319), .A3(113), .ZN(n396));
  INV_X1    g024(.A(322), .ZN(n397));
  NAND3_X1  g025(.A1(n397), .A2(319), .A3(101), .ZN(n398));
  INV_X1    g026(.A(319), .ZN(n399));
  NAND3_X1  g027(.A1(322), .A2(n399), .A3(125), .ZN(n400));
  NOR2_X1   g028(.A1(322), .A2(319), .ZN(n401));
  NAND2_X1  g029(.A1(n401), .A2(137), .ZN(n402));
  AND4_X1   g030(.A1(n400), .A2(n398), .A3(n396), .A4(n402), .ZN(1816));
  NAND3_X1  g031(.A1(322), .A2(319), .A3(112), .ZN(n404));
  NAND3_X1  g032(.A1(n397), .A2(319), .A3(100), .ZN(n405));
  NOR2_X1   g033(.A1(n397), .A2(319), .ZN(n406));
  AOI22_X1  g034(.A1(n406), .A2(124), .B1(136), .B2(n401), .ZN(n407));
  AND3_X1   g035(.A1(n407), .A2(n405), .A3(n404), .ZN(1817));
  AND3_X1   g036(.A1(322), .A2(319), .A3(114), .ZN(n409));
  AND3_X1   g037(.A1(n397), .A2(319), .A3(102), .ZN(n410));
  AND3_X1   g038(.A1(322), .A2(n399), .A3(126), .ZN(n411));
  AND2_X1   g039(.A1(n401), .A2(138), .ZN(n412));
  NOR4_X1   g040(.A1(n411), .A2(n410), .A3(n409), .A4(n412), .ZN(1818));
  NAND3_X1  g041(.A1(234), .A2(227), .A3(75), .ZN(n414));
  INV_X1    g042(.A(234), .ZN(n415));
  NAND3_X1  g043(.A1(n415), .A2(227), .A3(50), .ZN(n416));
  NOR2_X1   g044(.A1(n415), .A2(227), .ZN(n417));
  NOR2_X1   g045(.A1(234), .A2(227), .ZN(n418));
  AOI22_X1  g046(.A1(n417), .A2(62), .B1(88), .B2(n418), .ZN(n419));
  AND3_X1   g047(.A1(n419), .A2(n416), .A3(n414), .ZN(1819));
  AND2_X1   g048(.A1(n415), .A2(227), .ZN(n421));
  AND3_X1   g049(.A1(234), .A2(227), .A3(76), .ZN(n422));
  AOI21_X1  g050(.A(n422), .B1(n421), .B2(51), .ZN(n423));
  AOI22_X1  g051(.A1(n417), .A2(63), .B1(89), .B2(n418), .ZN(n424));
  NAND2_X1  g052(.A1(n424), .A2(n423), .ZN(2014));
  INV_X1    g053(.A(2014), .ZN(1820));
  NAND3_X1  g054(.A1(234), .A2(227), .A3(77), .ZN(n427));
  NAND3_X1  g055(.A1(n415), .A2(227), .A3(52), .ZN(n428));
  AOI22_X1  g056(.A1(n417), .A2(64), .B1(90), .B2(n418), .ZN(n429));
  AND3_X1   g057(.A1(n429), .A2(n428), .A3(n427), .ZN(1821));
  NAND3_X1  g058(.A1(234), .A2(227), .A3(68), .ZN(n431));
  NAND3_X1  g059(.A1(n415), .A2(227), .A3(43), .ZN(n432));
  AOI22_X1  g060(.A1(n417), .A2(56), .B1(81), .B2(n418), .ZN(n433));
  NAND4_X1  g061(.A1(n432), .A2(n431), .A3(241), .A4(n433), .ZN(1969));
  AND2_X1   g062(.A1(237), .A2(224), .ZN(n435));
  NAND3_X1  g063(.A1(n435), .A2(1726), .A3(36), .ZN(1970));
  NAND2_X1  g064(.A1(3), .A2(\1 ), .ZN(n437));
  NAND3_X1  g065(.A1(n437), .A2(n435), .A3(1726), .ZN(1971));
  NAND3_X1  g066(.A1(234), .A2(227), .A3(78), .ZN(n439));
  NAND3_X1  g067(.A1(n415), .A2(227), .A3(53), .ZN(n440));
  AOI22_X1  g068(.A1(n417), .A2(65), .B1(91), .B2(n418), .ZN(n441));
  NAND3_X1  g069(.A1(n441), .A2(n440), .A3(n439), .ZN(2010));
  INV_X1    g070(.A(1821), .ZN(2012));
  INV_X1    g071(.A(1819), .ZN(2016));
  INV_X1    g072(.A(74), .ZN(n445));
  AOI21_X1  g073(.A(n415), .B1(227), .B2(n445), .ZN(n446));
  AOI221_X1 g074(.A(n446), .B1(n421), .B2(49), .C1(87), .C2(n418), .ZN(n447));
  INV_X1    g075(.A(n447), .ZN(2018));
  NAND3_X1  g076(.A1(234), .A2(227), .A3(73), .ZN(n449));
  NAND3_X1  g077(.A1(n415), .A2(227), .A3(48), .ZN(n450));
  AOI22_X1  g078(.A1(n417), .A2(61), .B1(86), .B2(n418), .ZN(n451));
  AND3_X1   g079(.A1(n451), .A2(n450), .A3(n449), .ZN(n452));
  INV_X1    g080(.A(n452), .ZN(2020));
  NAND3_X1  g081(.A1(234), .A2(227), .A3(72), .ZN(n454));
  NAND3_X1  g082(.A1(n415), .A2(227), .A3(47), .ZN(n455));
  AOI22_X1  g083(.A1(n417), .A2(60), .B1(85), .B2(n418), .ZN(n456));
  AND3_X1   g084(.A1(n456), .A2(n455), .A3(n454), .ZN(n457));
  INV_X1    g085(.A(n457), .ZN(2022));
  INV_X1    g086(.A(246), .ZN(n459));
  NAND3_X1  g087(.A1(234), .A2(227), .A3(79), .ZN(n460));
  NAND3_X1  g088(.A1(n415), .A2(227), .A3(54), .ZN(n461));
  AOI22_X1  g089(.A1(n417), .A2(66), .B1(92), .B2(n418), .ZN(n462));
  AND3_X1   g090(.A1(n462), .A2(n461), .A3(n460), .ZN(n463));
  INV_X1    g091(.A(n463), .ZN(n464));
  MUX2_X1   g092(.S(n459), .B(n464), .A(2012), .Z(2387));
  MUX2_X1   g093(.S(n459), .B(2010), .A(2014), .Z(2389));
  INV_X1    g094(.A(230), .ZN(n467));
  OAI21_X1  g095(.A(n463), .B1(241), .B2(n467), .ZN(2496));
  AND3_X1   g096(.A1(n433), .A2(n432), .A3(n431), .ZN(n469));
  INV_X1    g097(.A(n469), .ZN(n470));
  AND4_X1   g098(.A1(n461), .A2(n460), .A3(n467), .A4(n462), .ZN(n471));
  INV_X1    g099(.A(n471), .ZN(n472));
  MUX2_X1   g100(.S(246), .B(n472), .A(n470), .Z(2643));
  NAND3_X1  g101(.A1(322), .A2(319), .A3(111), .ZN(n474));
  NAND3_X1  g102(.A1(n397), .A2(319), .A3(99), .ZN(n475));
  AOI22_X1  g103(.A1(n406), .A2(123), .B1(135), .B2(n401), .ZN(n476));
  AND3_X1   g104(.A1(n476), .A2(n475), .A3(n474), .ZN(n477));
  NOR2_X1   g105(.A1(n477), .A2(313), .ZN(n478));
  OR2_X1    g106(.A1(n478), .A2(n477), .ZN(n479));
  AND2_X1   g107(.A1(322), .A2(319), .ZN(n480));
  NOR2_X1   g108(.A1(322), .A2(n399), .ZN(n481));
  NOR4_X1   g109(.A1(n406), .A2(n481), .A3(n480), .A4(n401), .ZN(n482));
  XNOR2_X1  g110(.A(n482), .B(316), .ZN(n483));
  OAI211_X1 g111(.A(n479), .B(n483), .C1(n478), .C2(313), .ZN(2891));
  XOR2_X1   g112(.A(349), .B(346), .Z(n485));
  XNOR2_X1  g113(.A(259), .B(256), .ZN(n486));
  XNOR2_X1  g114(.A(n486), .B(n485), .ZN(n487));
  XNOR2_X1  g115(.A(331), .B(328), .ZN(n488));
  XNOR2_X1  g116(.A(343), .B(340), .ZN(n489));
  INV_X1    g117(.A(n489), .ZN(n490));
  XNOR2_X1  g118(.A(337), .B(334), .ZN(n491));
  INV_X1    g119(.A(n491), .ZN(n492));
  NOR3_X1   g120(.A1(n492), .A2(n490), .A3(n488), .ZN(n493));
  NOR3_X1   g121(.A1(n491), .A2(n489), .A3(n488), .ZN(n494));
  INV_X1    g122(.A(n488), .ZN(n495));
  NOR3_X1   g123(.A1(n492), .A2(n489), .A3(n495), .ZN(n496));
  NOR3_X1   g124(.A1(n491), .A2(n490), .A3(n495), .ZN(n497));
  NOR4_X1   g125(.A1(n496), .A2(n494), .A3(n493), .A4(n497), .ZN(n498));
  OAI21_X1  g126(.A(14), .B1(n498), .B2(n487), .ZN(n499));
  AOI21_X1  g127(.A(n499), .B1(n498), .B2(n487), .ZN(2925));
  XNOR2_X1  g128(.A(316), .B(313), .ZN(n501));
  XNOR2_X1  g129(.A(355), .B(294), .ZN(n502));
  XNOR2_X1  g130(.A(309), .B(305), .ZN(n503));
  INV_X1    g131(.A(n503), .ZN(n504));
  XNOR2_X1  g132(.A(301), .B(297), .ZN(n505));
  INV_X1    g133(.A(n505), .ZN(n506));
  NOR3_X1   g134(.A1(n506), .A2(n504), .A3(n502), .ZN(n507));
  NOR3_X1   g135(.A1(n505), .A2(n503), .A3(n502), .ZN(n508));
  INV_X1    g136(.A(n502), .ZN(n509));
  NOR3_X1   g137(.A1(n506), .A2(n503), .A3(n509), .ZN(n510));
  NOR3_X1   g138(.A1(n505), .A2(n504), .A3(n509), .ZN(n511));
  NOR4_X1   g139(.A1(n510), .A2(n508), .A3(n507), .A4(n511), .ZN(n512));
  XNOR2_X1  g140(.A(n512), .B(n501), .ZN(2970));
  XNOR2_X1  g141(.A(281), .B(278), .ZN(n514));
  XNOR2_X1  g142(.A(287), .B(284), .ZN(n515));
  XNOR2_X1  g143(.A(n515), .B(n514), .ZN(n516));
  XNOR2_X1  g144(.A(352), .B(263), .ZN(n517));
  XNOR2_X1  g145(.A(275), .B(272), .ZN(n518));
  INV_X1    g146(.A(n518), .ZN(n519));
  XNOR2_X1  g147(.A(269), .B(266), .ZN(n520));
  INV_X1    g148(.A(n520), .ZN(n521));
  NOR3_X1   g149(.A1(n521), .A2(n519), .A3(n517), .ZN(n522));
  NOR3_X1   g150(.A1(n520), .A2(n518), .A3(n517), .ZN(n523));
  INV_X1    g151(.A(n517), .ZN(n524));
  NOR3_X1   g152(.A1(n521), .A2(n518), .A3(n524), .ZN(n525));
  NOR3_X1   g153(.A1(n520), .A2(n519), .A3(n524), .ZN(n526));
  NOR4_X1   g154(.A1(n525), .A2(n523), .A3(n522), .A4(n526), .ZN(n527));
  XNOR2_X1  g155(.A(n527), .B(n516), .ZN(2971));
  MUX2_X1   g156(.S(16), .B(2014), .A(21), .Z(n529));
  MUX2_X1   g157(.S(16), .B(2016), .A(22), .Z(n530));
  XNOR2_X1  g158(.A(n530), .B(272), .ZN(n531));
  INV_X1    g159(.A(278), .ZN(n532));
  MUX2_X1   g160(.S(16), .B(2020), .A(6), .Z(n533));
  XNOR2_X1  g161(.A(n533), .B(n532), .ZN(n534));
  INV_X1    g162(.A(275), .ZN(n535));
  MUX2_X1   g163(.S(16), .B(2018), .A(23), .Z(n536));
  XNOR2_X1  g164(.A(n536), .B(n535), .ZN(n537));
  INV_X1    g165(.A(281), .ZN(n538));
  MUX2_X1   g166(.S(16), .B(2022), .A(24), .Z(n539));
  XNOR2_X1  g167(.A(n539), .B(n538), .ZN(n540));
  INV_X1    g168(.A(25), .ZN(n541));
  NAND3_X1  g169(.A1(322), .A2(319), .A3(107), .ZN(n542));
  NAND3_X1  g170(.A1(n397), .A2(319), .A3(95), .ZN(n543));
  AOI22_X1  g171(.A1(n406), .A2(119), .B1(131), .B2(n401), .ZN(n544));
  AND3_X1   g172(.A1(n544), .A2(n543), .A3(n542), .ZN(n545));
  MUX2_X1   g173(.S(29), .B(n545), .A(n541), .Z(n546));
  XNOR2_X1  g174(.A(n546), .B(284), .ZN(n547));
  NAND4_X1  g175(.A1(n540), .A2(n537), .A3(n534), .A4(n547), .ZN(n548));
  AOI211_X1 g176(.A(n531), .B(n548), .C1(n529), .C2(269), .ZN(n549));
  INV_X1    g177(.A(305), .ZN(n550));
  INV_X1    g178(.A(34), .ZN(n551));
  MUX2_X1   g179(.S(29), .B(1816), .A(n551), .Z(n552));
  NAND2_X1  g180(.A1(n459), .A2(11), .ZN(n553));
  NAND2_X1  g181(.A1(246), .A2(11), .ZN(n554));
  INV_X1    g182(.A(28), .ZN(n555));
  MUX2_X1   g183(.S(29), .B(n477), .A(n555), .Z(n556));
  AOI221_X1 g184(.A(n556), .B1(n553), .B2(n554), .C1(n552), .C2(n550), .ZN(n557));
  INV_X1    g185(.A(294), .ZN(n558));
  NAND3_X1  g186(.A1(322), .A2(319), .A3(115), .ZN(n559));
  NAND3_X1  g187(.A1(n397), .A2(319), .A3(103), .ZN(n560));
  AOI22_X1  g188(.A1(n406), .A2(127), .B1(139), .B2(n401), .ZN(n561));
  AND3_X1   g189(.A1(n561), .A2(n560), .A3(n559), .ZN(n562));
  INV_X1    g190(.A(n562), .ZN(n563));
  MUX2_X1   g191(.S(29), .B(n563), .A(33), .Z(n564));
  OAI22_X1  g192(.A1(n552), .A2(n550), .B1(297), .B2(n564), .ZN(n565));
  INV_X1    g193(.A(26), .ZN(n566));
  NAND3_X1  g194(.A1(322), .A2(319), .A3(116), .ZN(n567));
  NAND3_X1  g195(.A1(n397), .A2(319), .A3(104), .ZN(n568));
  AOI22_X1  g196(.A1(n406), .A2(128), .B1(140), .B2(n401), .ZN(n569));
  AND3_X1   g197(.A1(n569), .A2(n568), .A3(n567), .ZN(n570));
  MUX2_X1   g198(.S(29), .B(n570), .A(n566), .Z(n571));
  AOI221_X1 g199(.A(n565), .B1(n564), .B2(297), .C1(n558), .C2(n571), .ZN(n572));
  INV_X1    g200(.A(309), .ZN(n573));
  INV_X1    g201(.A(35), .ZN(n574));
  MUX2_X1   g202(.S(29), .B(1817), .A(n574), .Z(n575));
  NOR2_X1   g203(.A1(n575), .A2(n573), .ZN(n576));
  OR4_X1    g204(.A1(n411), .A2(n410), .A3(n409), .A4(n412), .ZN(n577));
  MUX2_X1   g205(.S(29), .B(n577), .A(27), .Z(n578));
  MUX2_X1   g206(.S(16), .B(2012), .A(5), .Z(n579));
  XNOR2_X1  g207(.A(n579), .B(266), .ZN(n580));
  AOI211_X1 g208(.A(n576), .B(n580), .C1(n578), .C2(301), .ZN(n581));
  NAND3_X1  g209(.A1(322), .A2(319), .A3(117), .ZN(n582));
  NAND3_X1  g210(.A1(n397), .A2(319), .A3(105), .ZN(n583));
  AOI22_X1  g211(.A1(n406), .A2(129), .B1(141), .B2(n401), .ZN(n584));
  NAND3_X1  g212(.A1(n584), .A2(n583), .A3(n582), .ZN(n585));
  MUX2_X1   g213(.S(29), .B(n585), .A(32), .Z(n586));
  OAI22_X1  g214(.A1(n571), .A2(n558), .B1(287), .B2(n586), .ZN(n587));
  AOI221_X1 g215(.A(n587), .B1(n575), .B2(n573), .C1(287), .C2(n586), .ZN(n588));
  MUX2_X1   g216(.S(16), .B(n464), .A(4), .Z(n589));
  XNOR2_X1  g217(.A(n589), .B(259), .ZN(n590));
  MUX2_X1   g218(.S(16), .B(n470), .A(19), .Z(n591));
  XNOR2_X1  g219(.A(n591), .B(256), .ZN(n592));
  OAI22_X1  g220(.A1(n529), .A2(269), .B1(301), .B2(n578), .ZN(n593));
  MUX2_X1   g221(.S(16), .B(2010), .A(20), .Z(n594));
  XNOR2_X1  g222(.A(n594), .B(263), .ZN(n595));
  NOR4_X1   g223(.A1(n593), .A2(n592), .A3(n590), .A4(n595), .ZN(n596));
  AND3_X1   g224(.A1(n596), .A2(n588), .A3(n581), .ZN(n597));
  AND4_X1   g225(.A1(n572), .A2(n557), .A3(n549), .A4(n597), .ZN(3038));
  NAND4_X1  g226(.A1(n572), .A2(n557), .A3(n549), .A4(n597), .ZN(3079));
  NAND3_X1  g227(.A1(234), .A2(227), .A3(80), .ZN(n600));
  NAND3_X1  g228(.A1(n415), .A2(227), .A3(55), .ZN(n601));
  AOI22_X1  g229(.A1(n417), .A2(67), .B1(93), .B2(n418), .ZN(n602));
  AND3_X1   g230(.A1(n602), .A2(n601), .A3(n600), .ZN(n603));
  INV_X1    g231(.A(n603), .ZN(n604));
  XNOR2_X1  g232(.A(n463), .B(n469), .ZN(n605));
  XNOR2_X1  g233(.A(n605), .B(n471), .ZN(n606));
  XNOR2_X1  g234(.A(n603), .B(n606), .ZN(n607));
  MUX2_X1   g235(.S(241), .B(n604), .A(n607), .Z(3546));
  XOR2_X1   g236(.A(1817), .B(1816), .Z(n609));
  XNOR2_X1  g237(.A(n482), .B(n477), .ZN(n610));
  XNOR2_X1  g238(.A(n610), .B(n609), .ZN(n611));
  NAND3_X1  g239(.A1(322), .A2(319), .A3(118), .ZN(n612));
  NAND3_X1  g240(.A1(n397), .A2(319), .A3(106), .ZN(n613));
  AOI22_X1  g241(.A1(n406), .A2(130), .B1(142), .B2(n401), .ZN(n614));
  AND3_X1   g242(.A1(n614), .A2(n613), .A3(n612), .ZN(n615));
  XNOR2_X1  g243(.A(n615), .B(n545), .ZN(n616));
  XNOR2_X1  g244(.A(n562), .B(n577), .ZN(n617));
  AND3_X1   g245(.A1(n584), .A2(n583), .A3(n582), .ZN(n618));
  XOR2_X1   g246(.A(n618), .B(n570), .Z(n619));
  NOR3_X1   g247(.A1(n619), .A2(n617), .A3(n616), .ZN(n620));
  XOR2_X1   g248(.A(n562), .B(n577), .Z(n621));
  XNOR2_X1  g249(.A(n618), .B(n570), .ZN(n622));
  NOR3_X1   g250(.A1(n622), .A2(n621), .A3(n616), .ZN(n623));
  XOR2_X1   g251(.A(n615), .B(n545), .Z(n624));
  NOR3_X1   g252(.A1(n619), .A2(n621), .A3(n624), .ZN(n625));
  NOR3_X1   g253(.A1(n622), .A2(n617), .A3(n624), .ZN(n626));
  NOR4_X1   g254(.A1(n625), .A2(n623), .A3(n620), .A4(n626), .ZN(n627));
  INV_X1    g255(.A(37), .ZN(n628));
  OAI21_X1  g256(.A(n628), .B1(n627), .B2(n611), .ZN(n629));
  AOI21_X1  g257(.A(n629), .B1(n627), .B2(n611), .ZN(3671));
  XOR2_X1   g258(.A(n447), .B(1819), .Z(n631));
  XNOR2_X1  g259(.A(n457), .B(n452), .ZN(n632));
  XNOR2_X1  g260(.A(n632), .B(n631), .ZN(n633));
  XOR2_X1   g261(.A(n603), .B(n469), .Z(n634));
  XNOR2_X1  g262(.A(n463), .B(2010), .ZN(n635));
  NOR3_X1   g263(.A1(n635), .A2(n634), .A3(n471), .ZN(n636));
  XNOR2_X1  g264(.A(n603), .B(n469), .ZN(n637));
  XOR2_X1   g265(.A(n463), .B(2010), .Z(n638));
  NOR3_X1   g266(.A1(n638), .A2(n637), .A3(n471), .ZN(n639));
  NOR3_X1   g267(.A1(n638), .A2(n634), .A3(n472), .ZN(n640));
  NOR3_X1   g268(.A1(n635), .A2(n637), .A3(n472), .ZN(n641));
  NOR4_X1   g269(.A1(n640), .A2(n639), .A3(n636), .A4(n641), .ZN(n642));
  XNOR2_X1  g270(.A(n642), .B(n633), .ZN(n643));
  MUX2_X1   g271(.S(246), .B(n643), .A(n604), .Z(3803));
  XNOR2_X1  g272(.A(1821), .B(2014), .ZN(n645));
  NOR3_X1   g273(.A1(n645), .A2(n635), .A3(n637), .ZN(n646));
  XOR2_X1   g274(.A(1821), .B(2014), .Z(n647));
  NOR3_X1   g275(.A1(n647), .A2(n638), .A3(n637), .ZN(n648));
  NOR3_X1   g276(.A1(n647), .A2(n635), .A3(n634), .ZN(n649));
  NOR3_X1   g277(.A1(n645), .A2(n638), .A3(n634), .ZN(n650));
  NOR4_X1   g278(.A1(n649), .A2(n648), .A3(n646), .A4(n650), .ZN(n651));
  OAI21_X1  g279(.A(n628), .B1(n651), .B2(n633), .ZN(n652));
  AOI21_X1  g280(.A(n652), .B1(n651), .B2(n633), .ZN(3809));
  INV_X1    g281(.A(40), .ZN(n654));
  NAND4_X1  g282(.A1(n400), .A2(n398), .A3(n396), .A4(n402), .ZN(n655));
  NOR4_X1   g283(.A1(n655), .A2(262), .A3(n654), .A4(1818), .ZN(n656));
  OAI211_X1 g284(.A(1816), .B(40), .C1(262), .C2(1818), .ZN(n657));
  OR3_X1    g285(.A1(n657), .A2(n656), .A3(294), .ZN(n658));
  NOR3_X1   g286(.A1(n657), .A2(n656), .A3(n570), .ZN(n659));
  XNOR2_X1  g287(.A(n659), .B(n658), .ZN(n660));
  OR3_X1    g288(.A1(n657), .A2(n656), .A3(287), .ZN(n661));
  NOR3_X1   g289(.A1(n657), .A2(n656), .A3(n618), .ZN(n662));
  XNOR2_X1  g290(.A(n662), .B(n661), .ZN(n663));
  OR3_X1    g291(.A1(n657), .A2(n656), .A3(284), .ZN(n664));
  NOR3_X1   g292(.A1(n657), .A2(n656), .A3(n545), .ZN(n665));
  NOR4_X1   g293(.A1(n664), .A2(n663), .A3(n660), .A4(n665), .ZN(n666));
  INV_X1    g294(.A(262), .ZN(n667));
  NAND4_X1  g295(.A1(1816), .A2(n667), .A3(40), .A4(n577), .ZN(n668));
  INV_X1    g296(.A(n657), .ZN(n669));
  NAND4_X1  g297(.A1(n668), .A2(n457), .A3(n538), .A4(n669), .ZN(n670));
  XNOR2_X1  g298(.A(n665), .B(n664), .ZN(n671));
  NOR4_X1   g299(.A1(n670), .A2(n663), .A3(n660), .A4(n671), .ZN(n672));
  OR2_X1    g300(.A1(n659), .A2(n658), .ZN(n673));
  OR4_X1    g301(.A1(n656), .A2(n585), .A3(287), .A4(n657), .ZN(n674));
  OAI21_X1  g302(.A(n673), .B1(n674), .B2(n660), .ZN(n675));
  NOR3_X1   g303(.A1(n675), .A2(n672), .A3(n666), .ZN(n676));
  MUX2_X1   g304(.S(n656), .B(297), .A(263), .Z(n677));
  XOR2_X1   g305(.A(n677), .B(2010), .Z(n678));
  INV_X1    g306(.A(259), .ZN(n679));
  MUX2_X1   g307(.S(n668), .B(n679), .A(n558), .Z(n680));
  XNOR2_X1  g308(.A(n680), .B(n464), .ZN(n681));
  OR2_X1    g309(.A1(n668), .A2(287), .ZN(n682));
  OAI21_X1  g310(.A(n682), .B1(n656), .B2(256), .ZN(n683));
  NAND4_X1  g311(.A1(n681), .A2(n678), .A3(n469), .A4(n683), .ZN(n684));
  NAND3_X1  g312(.A1(n680), .A2(n678), .A3(n463), .ZN(n685));
  OAI211_X1 g313(.A(n684), .B(n685), .C1(n677), .C2(2010), .ZN(n686));
  INV_X1    g314(.A(8), .ZN(n687));
  MUX2_X1   g315(.S(n656), .B(309), .A(272), .Z(n688));
  NOR2_X1   g316(.A1(n688), .A2(n687), .ZN(n689));
  OR2_X1    g317(.A1(1819), .A2(n687), .ZN(n690));
  XNOR2_X1  g318(.A(n690), .B(n689), .ZN(n691));
  MUX2_X1   g319(.S(n656), .B(305), .A(269), .Z(n692));
  NOR2_X1   g320(.A1(n692), .A2(n687), .ZN(n693));
  NAND2_X1  g321(.A1(2014), .A2(8), .ZN(n694));
  XNOR2_X1  g322(.A(n694), .B(n693), .ZN(n695));
  MUX2_X1   g323(.S(n656), .B(301), .A(266), .Z(n696));
  XNOR2_X1  g324(.A(n696), .B(1821), .ZN(n697));
  NOR3_X1   g325(.A1(n656), .A2(275), .A3(n687), .ZN(n698));
  NOR3_X1   g326(.A1(n656), .A2(n447), .A3(n687), .ZN(n699));
  XNOR2_X1  g327(.A(n699), .B(n698), .ZN(n700));
  NOR3_X1   g328(.A1(n656), .A2(278), .A3(n687), .ZN(n701));
  NOR3_X1   g329(.A1(n656), .A2(n452), .A3(n687), .ZN(n702));
  XNOR2_X1  g330(.A(n702), .B(n701), .ZN(n703));
  NAND3_X1  g331(.A1(n703), .A2(n700), .A3(n697), .ZN(n704));
  NOR3_X1   g332(.A1(n704), .A2(n695), .A3(n691), .ZN(n705));
  NOR2_X1   g333(.A1(n696), .A2(2012), .ZN(n706));
  NAND3_X1  g334(.A1(n706), .A2(n703), .A3(n700), .ZN(n707));
  NOR3_X1   g335(.A1(n707), .A2(n695), .A3(n691), .ZN(n708));
  NAND4_X1  g336(.A1(n700), .A2(n694), .A3(n693), .A4(n703), .ZN(n709));
  NAND4_X1  g337(.A1(n700), .A2(n690), .A3(n689), .A4(n703), .ZN(n710));
  AND4_X1   g338(.A1(n452), .A2(n532), .A3(8), .A4(n668), .ZN(n711));
  AND4_X1   g339(.A1(n447), .A2(n535), .A3(8), .A4(n668), .ZN(n712));
  AOI21_X1  g340(.A(n711), .B1(n712), .B2(n703), .ZN(n713));
  OAI211_X1 g341(.A(n710), .B(n713), .C1(n709), .C2(n691), .ZN(n714));
  AOI211_X1 g342(.A(n708), .B(n714), .C1(n705), .C2(n686), .ZN(n715));
  NOR3_X1   g343(.A1(n657), .A2(n656), .A3(n457), .ZN(n716));
  NOR3_X1   g344(.A1(n657), .A2(n656), .A3(281), .ZN(n717));
  XOR2_X1   g345(.A(n717), .B(n716), .Z(n718));
  OR4_X1    g346(.A1(n671), .A2(n663), .A3(n660), .A4(n718), .ZN(n719));
  OAI21_X1  g347(.A(n676), .B1(n719), .B2(n715), .ZN(3851));
  LOGIC0_X1 g348(.Z(3875));
  INV_X1    g349(.A(1726), .ZN(n722));
  OR4_X1    g350(.A1(2970), .A2(2925), .A3(n722), .A4(2971), .ZN(n723));
  NOR3_X1   g351(.A1(n723), .A2(3809), .A3(3671), .ZN(3881));
  OR3_X1    g352(.A1(n723), .A2(3809), .A3(3671), .ZN(3882));
  BUF_X1    g353(.A(219), .Z(398));
  BUF_X1    g354(.A(219), .Z(400));
  BUF_X1    g355(.A(219), .Z(401));
  BUF_X1    g356(.A(253), .Z(419));
  BUF_X1    g357(.A(253), .Z(420));
  BUF_X1    g358(.A(290), .Z(456));
  BUF_X1    g359(.A(290), .Z(457));
  BUF_X1    g360(.A(290), .Z(458));
  BUF_X1    g361(.A(219), .Z(805));
  MUX2_X1   g362(.S(n459), .B(n464), .A(2012), .Z(2388));
  MUX2_X1   g363(.S(n459), .B(2010), .A(2014), .Z(2390));
  MUX2_X1   g364(.S(246), .B(n472), .A(n470), .Z(2644));
  MUX2_X1   g365(.S(246), .B(n643), .A(n604), .Z(3804));
endmodule


