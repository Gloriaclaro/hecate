// Benchmark "c1908" written by ABC on Tue Dec 06 12:35:31 2022

module c1908 ( 
    \1 , 4, 7, 10, 13, 16, 19, 22, 25, 28, 31, 34, 37, 40, 43, 46, 49, 53,
    56, 60, 63, 66, 69, 72, 76, 79, 82, 85, 88, 91, 94, 99, 104,
    2753, 2754, 2755, 2756, 2762, 2767, 2768, 2779, 2780, 2781, 2782, 2783,
    2784, 2785, 2786, 2787, 2811, 2886, 2887, 2888, 2889, 2890, 2891, 2892,
    2899  );
  input  \1 , 4, 7, 10, 13, 16, 19, 22, 25, 28, 31, 34, 37, 40, 43, 46,
    49, 53, 56, 60, 63, 66, 69, 72, 76, 79, 82, 85, 88, 91, 94, 99, 104;
  output 2753, 2754, 2755, 2756, 2762, 2767, 2768, 2779, 2780, 2781, 2782,
    2783, 2784, 2785, 2786, 2787, 2811, 2886, 2887, 2888, 2889, 2890, 2891,
    2892, 2899;
  wire n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
    n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
    n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
    n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
    n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
    n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
    n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
    n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n159, n160,
    n161, n162, n163, n164, n165, n166, n167, n168, n170, n171, n173, n174,
    n175, n176, n177, n179, n180, n181, n182, n183, n184, n186, n187, n188,
    n189, n190, n192, n193, n195, n196, n197, n198, n200, n202, n203, n204,
    n206, n207, n208, n210, n211, n213, n214, n215, n217, n219, n220, n221,
    n223, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
    n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
    n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
    n260, n262, n263, n264, n266, n267, n269, n270, n271, n273, n274, n276,
    n277, n279, n280, n281, n282, n284, n285, n286, n287, n288, n289, n290,
    n292, n293, n294;
  INV_X1    g000(.A(\1 ), .ZN(n58));
  INV_X1    g001(.A(94), .ZN(n59));
  INV_X1    g002(.A(46), .ZN(n60));
  XNOR2_X1  g003(.A(40), .B(25), .ZN(n61));
  XNOR2_X1  g004(.A(n61), .B(n60), .ZN(n62));
  XNOR2_X1  g005(.A(28), .B(19), .ZN(n63));
  XNOR2_X1  g006(.A(n63), .B(10), .ZN(n64));
  XNOR2_X1  g007(.A(n64), .B(n62), .ZN(n65));
  INV_X1    g008(.A(37), .ZN(n66));
  INV_X1    g009(.A(60), .ZN(n67));
  INV_X1    g010(.A(69), .ZN(n68));
  NOR3_X1   g011(.A1(104), .A2(n68), .A3(n67), .ZN(n69));
  XNOR2_X1  g012(.A(n69), .B(n66), .ZN(n70));
  XOR2_X1   g013(.A(n70), .B(n65), .Z(n71));
  AND2_X1   g014(.A1(n71), .A2(n59), .ZN(n72));
  INV_X1    g015(.A(56), .ZN(n73));
  AOI21_X1  g016(.A(n73), .B1(n59), .B2(69), .ZN(n74));
  INV_X1    g017(.A(n74), .ZN(n75));
  XNOR2_X1  g018(.A(n75), .B(n72), .ZN(n76));
  INV_X1    g019(.A(49), .ZN(n77));
  OR2_X1    g020(.A1(104), .A2(72), .ZN(n78));
  NOR2_X1   g021(.A1(n78), .A2(n77), .ZN(n79));
  XNOR2_X1  g022(.A(n79), .B(n58), .ZN(n80));
  INV_X1    g023(.A(13), .ZN(n81));
  XNOR2_X1  g024(.A(19), .B(16), .ZN(n82));
  XNOR2_X1  g025(.A(n82), .B(n81), .ZN(n83));
  XNOR2_X1  g026(.A(46), .B(43), .ZN(n84));
  XNOR2_X1  g027(.A(n84), .B(28), .ZN(n85));
  XNOR2_X1  g028(.A(37), .B(34), .ZN(n86));
  XNOR2_X1  g029(.A(n86), .B(31), .ZN(n87));
  XOR2_X1   g030(.A(n87), .B(n85), .Z(n88));
  XNOR2_X1  g031(.A(n88), .B(n83), .ZN(n89));
  XNOR2_X1  g032(.A(n89), .B(n80), .ZN(n90));
  OAI21_X1  g033(.A(79), .B1(n90), .B2(94), .ZN(n91));
  OR3_X1    g034(.A1(n90), .A2(94), .A3(79), .ZN(n92));
  AOI21_X1  g035(.A(n76), .B1(n92), .B2(n91), .ZN(n93));
  INV_X1    g036(.A(53), .ZN(n94));
  INV_X1    g037(.A(72), .ZN(n95));
  AOI21_X1  g038(.A(n94), .B1(n59), .B2(n95), .ZN(n96));
  INV_X1    g039(.A(n96), .ZN(n97));
  INV_X1    g040(.A(25), .ZN(n98));
  XNOR2_X1  g041(.A(n85), .B(n98), .ZN(n99));
  INV_X1    g042(.A(104), .ZN(n100));
  AND2_X1   g043(.A1(n100), .A2(63), .ZN(n101));
  XNOR2_X1  g044(.A(n101), .B(n99), .ZN(n102));
  XNOR2_X1  g045(.A(7), .B(4), .ZN(n103));
  XNOR2_X1  g046(.A(n103), .B(\1 ), .ZN(n104));
  XOR2_X1   g047(.A(n104), .B(n83), .Z(n105));
  XNOR2_X1  g048(.A(22), .B(10), .ZN(n106));
  XNOR2_X1  g049(.A(n106), .B(n105), .ZN(n107));
  OAI21_X1  g050(.A(n59), .B1(n107), .B2(n102), .ZN(n108));
  AOI21_X1  g051(.A(n108), .B1(n107), .B2(n102), .ZN(n109));
  AOI21_X1  g052(.A(n77), .B1(n59), .B2(n95), .ZN(n110));
  INV_X1    g053(.A(n110), .ZN(n111));
  XNOR2_X1  g054(.A(n111), .B(n109), .ZN(n112));
  AOI21_X1  g055(.A(n67), .B1(n59), .B2(69), .ZN(n113));
  XOR2_X1   g056(.A(40), .B(10), .Z(n114));
  AND2_X1   g057(.A1(n100), .A2(66), .ZN(n115));
  XOR2_X1   g058(.A(n115), .B(n114), .Z(n116));
  XNOR2_X1  g059(.A(n104), .B(n85), .ZN(n117));
  XNOR2_X1  g060(.A(n117), .B(n87), .ZN(n118));
  XNOR2_X1  g061(.A(n118), .B(n116), .ZN(n119));
  OAI21_X1  g062(.A(76), .B1(n119), .B2(94), .ZN(n120));
  INV_X1    g063(.A(76), .ZN(n121));
  XOR2_X1   g064(.A(n118), .B(n116), .Z(n122));
  NAND3_X1  g065(.A1(n122), .A2(n59), .A3(n121), .ZN(n123));
  AOI21_X1  g066(.A(n113), .B1(n123), .B2(n120), .ZN(n124));
  NAND4_X1  g067(.A1(n112), .A2(n97), .A3(n93), .A4(n124), .ZN(n125));
  AND2_X1   g068(.A1(72), .A2(69), .ZN(n126));
  NOR4_X1   g069(.A1(n100), .A2(n59), .A3(88), .A4(n126), .ZN(n127));
  INV_X1    g070(.A(99), .ZN(n128));
  NOR3_X1   g071(.A1(n126), .A2(104), .A3(n128), .ZN(n129));
  NOR2_X1   g072(.A1(n129), .A2(n127), .ZN(n130));
  INV_X1    g073(.A(n130), .ZN(n131));
  INV_X1    g074(.A(7), .ZN(n132));
  XNOR2_X1  g075(.A(22), .B(16), .ZN(n133));
  XNOR2_X1  g076(.A(n133), .B(n132), .ZN(n134));
  XNOR2_X1  g077(.A(43), .B(28), .ZN(n135));
  XNOR2_X1  g078(.A(n135), .B(34), .ZN(n136));
  XNOR2_X1  g079(.A(n136), .B(n134), .ZN(n137));
  NOR3_X1   g080(.A1(104), .A2(n68), .A3(n73), .ZN(n138));
  XNOR2_X1  g081(.A(n138), .B(n137), .ZN(n139));
  NOR2_X1   g082(.A1(n139), .A2(94), .ZN(n140));
  XNOR2_X1  g083(.A(n140), .B(85), .ZN(n141));
  NOR2_X1   g084(.A1(104), .A2(72), .ZN(n142));
  AOI21_X1  g085(.A(43), .B1(n142), .B2(53), .ZN(n143));
  INV_X1    g086(.A(43), .ZN(n144));
  NOR3_X1   g087(.A1(n78), .A2(n94), .A3(n144), .ZN(n145));
  OAI21_X1  g088(.A(31), .B1(n145), .B2(n143), .ZN(n146));
  OR3_X1    g089(.A1(n145), .A2(n143), .A3(31), .ZN(n147));
  AND3_X1   g090(.A1(n147), .A2(n146), .A3(n62), .ZN(n148));
  AOI21_X1  g091(.A(n62), .B1(n147), .B2(n146), .ZN(n149));
  XNOR2_X1  g092(.A(22), .B(13), .ZN(n150));
  XNOR2_X1  g093(.A(n150), .B(4), .ZN(n151));
  OAI21_X1  g094(.A(n151), .B1(n149), .B2(n148), .ZN(n152));
  OR3_X1    g095(.A1(n151), .A2(n149), .A3(n148), .ZN(n153));
  AOI21_X1  g096(.A(94), .B1(n153), .B2(n152), .ZN(n154));
  XNOR2_X1  g097(.A(n154), .B(82), .ZN(n155));
  NAND3_X1  g098(.A1(n155), .A2(n141), .A3(n131), .ZN(n156));
  NOR2_X1   g099(.A1(n156), .A2(n125), .ZN(n157));
  XNOR2_X1  g100(.A(n157), .B(n58), .ZN(2753));
  INV_X1    g101(.A(79), .ZN(n159));
  XOR2_X1   g102(.A(n89), .B(n80), .Z(n160));
  AOI21_X1  g103(.A(n159), .B1(n160), .B2(n59), .ZN(n161));
  NOR3_X1   g104(.A1(n90), .A2(94), .A3(79), .ZN(n162));
  NOR3_X1   g105(.A1(n162), .A2(n161), .A3(n76), .ZN(n163));
  NAND4_X1  g106(.A1(n124), .A2(n112), .A3(n97), .A4(n163), .ZN(n164));
  INV_X1    g107(.A(82), .ZN(n165));
  XNOR2_X1  g108(.A(n154), .B(n165), .ZN(n166));
  NAND3_X1  g109(.A1(n166), .A2(n141), .A3(n131), .ZN(n167));
  NOR2_X1   g110(.A1(n167), .A2(n164), .ZN(n168));
  XOR2_X1   g111(.A(n168), .B(4), .Z(2754));
  OR3_X1    g112(.A1(n166), .A2(n141), .A3(n130), .ZN(n170));
  NOR2_X1   g113(.A1(n170), .A2(n164), .ZN(n171));
  XNOR2_X1  g114(.A(n171), .B(n132), .ZN(2755));
  NAND3_X1  g115(.A1(n124), .A2(n112), .A3(n97), .ZN(n173));
  XNOR2_X1  g116(.A(n74), .B(n72), .ZN(n174));
  NOR3_X1   g117(.A1(n162), .A2(n161), .A3(n174), .ZN(n175));
  NAND4_X1  g118(.A1(n155), .A2(n141), .A3(n131), .A4(n175), .ZN(n176));
  NOR2_X1   g119(.A1(n176), .A2(n173), .ZN(n177));
  XOR2_X1   g120(.A(n177), .B(10), .Z(2756));
  AOI21_X1  g121(.A(n174), .B1(n92), .B2(n91), .ZN(n179));
  NAND4_X1  g122(.A1(n124), .A2(n112), .A3(n97), .A4(n179), .ZN(n180));
  NOR4_X1   g123(.A1(n100), .A2(n59), .A3(91), .A4(n126), .ZN(n181));
  NOR2_X1   g124(.A1(n181), .A2(n129), .ZN(n182));
  OR3_X1    g125(.A1(n182), .A2(n166), .A3(n141), .ZN(n183));
  OR2_X1    g126(.A1(n183), .A2(n180), .ZN(n184));
  XNOR2_X1  g127(.A(n184), .B(28), .ZN(2762));
  INV_X1    g128(.A(85), .ZN(n186));
  XNOR2_X1  g129(.A(n140), .B(n186), .ZN(n187));
  INV_X1    g130(.A(n182), .ZN(n188));
  NAND3_X1  g131(.A1(n188), .A2(n166), .A3(n187), .ZN(n189));
  NOR2_X1   g132(.A1(n189), .A2(n125), .ZN(n190));
  XNOR2_X1  g133(.A(n190), .B(n144), .ZN(2767));
  NAND3_X1  g134(.A1(n188), .A2(n166), .A3(n141), .ZN(n192));
  NOR2_X1   g135(.A1(n192), .A2(n180), .ZN(n193));
  XNOR2_X1  g136(.A(n193), .B(n60), .ZN(2768));
  INV_X1    g137(.A(n113), .ZN(n195));
  AND3_X1   g138(.A1(n123), .A2(n120), .A3(n195), .ZN(n196));
  NAND4_X1  g139(.A1(n112), .A2(n97), .A3(n93), .A4(n196), .ZN(n197));
  NOR2_X1   g140(.A1(n197), .A2(n167), .ZN(n198));
  XNOR2_X1  g141(.A(n198), .B(n81), .ZN(2779));
  NOR2_X1   g142(.A1(n197), .A2(n170), .ZN(n200));
  XOR2_X1   g143(.A(n200), .B(16), .Z(2780));
  NAND3_X1  g144(.A1(n196), .A2(n112), .A3(n97), .ZN(n202));
  NAND4_X1  g145(.A1(n155), .A2(n141), .A3(n131), .A4(n179), .ZN(n203));
  NOR2_X1   g146(.A1(n203), .A2(n202), .ZN(n204));
  XOR2_X1   g147(.A(n204), .B(19), .Z(2781));
  NAND4_X1  g148(.A1(n163), .A2(n112), .A3(n97), .A4(n196), .ZN(n206));
  NAND3_X1  g149(.A1(n166), .A2(n187), .A3(n131), .ZN(n207));
  NOR2_X1   g150(.A1(n207), .A2(n206), .ZN(n208));
  XOR2_X1   g151(.A(n208), .B(22), .Z(2782));
  NAND4_X1  g152(.A1(n175), .A2(n166), .A3(n141), .A4(n188), .ZN(n210));
  NOR2_X1   g153(.A1(n210), .A2(n202), .ZN(n211));
  XNOR2_X1  g154(.A(n211), .B(n98), .ZN(2783));
  XNOR2_X1  g155(.A(n110), .B(n109), .ZN(n213));
  NAND4_X1  g156(.A1(n213), .A2(n97), .A3(n93), .A4(n124), .ZN(n214));
  NOR2_X1   g157(.A1(n214), .A2(n192), .ZN(n215));
  XOR2_X1   g158(.A(n215), .B(31), .Z(2784));
  NOR2_X1   g159(.A1(n214), .A2(n183), .ZN(n217));
  XOR2_X1   g160(.A(n217), .B(34), .Z(2785));
  NAND3_X1  g161(.A1(n124), .A2(n213), .A3(n97), .ZN(n219));
  NAND4_X1  g162(.A1(n179), .A2(n155), .A3(n141), .A4(n188), .ZN(n220));
  NOR2_X1   g163(.A1(n220), .A2(n219), .ZN(n221));
  XNOR2_X1  g164(.A(n221), .B(n66), .ZN(2786));
  NOR2_X1   g165(.A1(n219), .A2(n210), .ZN(n223));
  XOR2_X1   g166(.A(n223), .B(40), .Z(2787));
  NAND4_X1  g167(.A1(n195), .A2(n97), .A3(n174), .A4(n141), .ZN(n225));
  NAND4_X1  g168(.A1(n120), .A2(n92), .A3(n91), .A4(n123), .ZN(n226));
  NOR4_X1   g169(.A1(n225), .A2(n166), .A3(n112), .A4(n226), .ZN(n227));
  NOR3_X1   g170(.A1(n227), .A2(104), .A3(99), .ZN(n228));
  OAI22_X1  g171(.A1(n176), .A2(n173), .B1(n167), .B2(n197), .ZN(n229));
  OAI22_X1  g172(.A1(n197), .A2(n170), .B1(n202), .B2(n203), .ZN(n230));
  OAI22_X1  g173(.A1(n206), .A2(n207), .B1(n167), .B2(n164), .ZN(n231));
  OAI22_X1  g174(.A1(n164), .A2(n170), .B1(n156), .B2(n125), .ZN(n232));
  NOR4_X1   g175(.A1(n231), .A2(n230), .A3(n229), .A4(n232), .ZN(n233));
  OAI22_X1  g176(.A1(n214), .A2(n183), .B1(n219), .B2(n220), .ZN(n234));
  OAI22_X1  g177(.A1(n210), .A2(n219), .B1(n189), .B2(n125), .ZN(n235));
  OAI22_X1  g178(.A1(n202), .A2(n210), .B1(n192), .B2(n180), .ZN(n236));
  OAI22_X1  g179(.A1(n192), .A2(n214), .B1(n183), .B2(n180), .ZN(n237));
  NOR4_X1   g180(.A1(n236), .A2(n235), .A3(n234), .A4(n237), .ZN(n238));
  AND2_X1   g181(.A1(n238), .A2(n233), .ZN(n239));
  AND3_X1   g182(.A1(n196), .A2(n213), .A3(n97), .ZN(n240));
  INV_X1    g183(.A(n129), .ZN(n241));
  NOR3_X1   g184(.A1(n166), .A2(n187), .A3(n241), .ZN(n242));
  NAND3_X1  g185(.A1(n242), .A2(n240), .A3(n93), .ZN(n243));
  NAND3_X1  g186(.A1(n242), .A2(n240), .A3(n175), .ZN(n244));
  NOR3_X1   g187(.A1(n166), .A2(n141), .A3(n241), .ZN(n245));
  NAND3_X1  g188(.A1(n245), .A2(n240), .A3(n163), .ZN(n246));
  NAND3_X1  g189(.A1(n246), .A2(n244), .A3(n243), .ZN(n247));
  NAND3_X1  g190(.A1(n163), .A2(n155), .A3(n141), .ZN(n248));
  NAND4_X1  g191(.A1(n129), .A2(n213), .A3(n96), .A4(n196), .ZN(n249));
  OR2_X1    g192(.A1(n248), .A2(n249), .ZN(n250));
  AND4_X1   g193(.A1(n123), .A2(n120), .A3(n113), .A4(n129), .ZN(n251));
  NAND3_X1  g194(.A1(n251), .A2(n213), .A3(n97), .ZN(n252));
  OAI211_X1 g195(.A(n250), .B(99), .C1(n248), .C2(n252), .ZN(n253));
  NAND3_X1  g196(.A1(n92), .A2(n91), .A3(n174), .ZN(n254));
  NAND3_X1  g197(.A1(n155), .A2(n141), .A3(n129), .ZN(n255));
  AOI211_X1 g198(.A(n254), .B(n255), .C1(n219), .C2(n202), .ZN(n256));
  NOR3_X1   g199(.A1(n155), .A2(n187), .A3(n241), .ZN(n257));
  AND3_X1   g200(.A1(n257), .A2(n240), .A3(n163), .ZN(n258));
  OR4_X1    g201(.A1(n256), .A2(n227), .A3(104), .A4(n258), .ZN(n259));
  NOR3_X1   g202(.A1(n259), .A2(n253), .A3(n247), .ZN(n260));
  AOI21_X1  g203(.A(n228), .B1(n260), .B2(n239), .ZN(2811));
  XOR2_X1   g204(.A(n107), .B(n102), .Z(n262));
  AOI211_X1 g205(.A(n111), .B(n59), .C1(n233), .C2(n238), .ZN(n263));
  XNOR2_X1  g206(.A(n263), .B(n262), .ZN(n264));
  AOI21_X1  g207(.A(n264), .B1(104), .B2(n128), .ZN(2886));
  AOI211_X1 g208(.A(n59), .B(n121), .C1(n233), .C2(n238), .ZN(n266));
  XNOR2_X1  g209(.A(n266), .B(n122), .ZN(n267));
  AOI21_X1  g210(.A(n267), .B1(104), .B2(n128), .ZN(2887));
  NAND2_X1  g211(.A1(n153), .A2(n152), .ZN(n269));
  AOI211_X1 g212(.A(n59), .B(n165), .C1(n233), .C2(n238), .ZN(n270));
  XNOR2_X1  g213(.A(n270), .B(n269), .ZN(n271));
  AOI21_X1  g214(.A(n271), .B1(104), .B2(n128), .ZN(2888));
  AOI211_X1 g215(.A(n59), .B(n186), .C1(n233), .C2(n238), .ZN(n273));
  XOR2_X1   g216(.A(n273), .B(n139), .Z(n274));
  AOI21_X1  g217(.A(n274), .B1(104), .B2(n128), .ZN(2889));
  AOI211_X1 g218(.A(n75), .B(n59), .C1(n233), .C2(n238), .ZN(n276));
  XNOR2_X1  g219(.A(n276), .B(n71), .ZN(n277));
  AOI21_X1  g220(.A(n277), .B1(104), .B2(n128), .ZN(2890));
  OR2_X1    g221(.A1(n233), .A2(104), .ZN(n279));
  OAI21_X1  g222(.A(n107), .B1(n100), .B2(88), .ZN(n280));
  XNOR2_X1  g223(.A(n280), .B(n279), .ZN(n281));
  AOI21_X1  g224(.A(n100), .B1(88), .B2(63), .ZN(n282));
  XNOR2_X1  g225(.A(n282), .B(n281), .ZN(2891));
  NOR2_X1   g226(.A1(n238), .A2(104), .ZN(n284));
  OR2_X1    g227(.A1(n88), .A2(n61), .ZN(n285));
  NOR2_X1   g228(.A1(n100), .A2(91), .ZN(n286));
  AOI21_X1  g229(.A(n286), .B1(n88), .B2(n61), .ZN(n287));
  AND2_X1   g230(.A1(n287), .A2(n285), .ZN(n288));
  XNOR2_X1  g231(.A(n288), .B(n284), .ZN(n289));
  AOI21_X1  g232(.A(n100), .B1(91), .B2(66), .ZN(n290));
  XNOR2_X1  g233(.A(n290), .B(n289), .ZN(2892));
  AOI211_X1 g234(.A(n59), .B(n159), .C1(n233), .C2(n238), .ZN(n292));
  XOR2_X1   g235(.A(n292), .B(n89), .Z(n293));
  XNOR2_X1  g236(.A(n293), .B(n80), .ZN(n294));
  AOI21_X1  g237(.A(n294), .B1(104), .B2(n128), .ZN(2899));
endmodule


