// Benchmark "c499" written by ABC on Tue Dec 06 12:34:27 2022

module c499 ( 
    \1 , 5, 9, 13, 17, 21, 25, 29, 33, 37, 41, 45, 49, 53, 57, 61, 65, 69,
    73, 77, 81, 85, 89, 93, 97, 101, 105, 109, 113, 117, 121, 125, 129,
    130, 131, 132, 133, 134, 135, 136, 137,
    724, 725, 726, 727, 728, 729, 730, 731, 732, 733, 734, 735, 736, 737,
    738, 739, 740, 741, 742, 743, 744, 745, 746, 747, 748, 749, 750, 751,
    752, 753, 754, 755  );
  input  \1 , 5, 9, 13, 17, 21, 25, 29, 33, 37, 41, 45, 49, 53, 57, 61,
    65, 69, 73, 77, 81, 85, 89, 93, 97, 101, 105, 109, 113, 117, 121, 125,
    129, 130, 131, 132, 133, 134, 135, 136, 137;
  output 724, 725, 726, 727, 728, 729, 730, 731, 732, 733, 734, 735, 736, 737,
    738, 739, 740, 741, 742, 743, 744, 745, 746, 747, 748, 749, 750, 751,
    752, 753, 754, 755;
  wire n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
    n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
    n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
    n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
    n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
    n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
    n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
    n161, n162, n163, n164, n166, n168, n170, n172, n173, n174, n176, n178,
    n180, n182, n183, n184, n185, n187, n189, n191, n193, n194, n196, n198,
    n200, n202, n203, n204, n205, n206, n207, n208, n209, n210, n212, n214,
    n216, n218, n219, n221, n223, n225, n227, n228, n230, n232, n234, n236,
    n237, n239, n241, n243;
  XNOR2_X1  g000(.A(17), .B(\1 ), .ZN(n73));
  XNOR2_X1  g001(.A(49), .B(33), .ZN(n74));
  XNOR2_X1  g002(.A(n74), .B(n73), .ZN(n75));
  NAND2_X1  g003(.A1(137), .A2(129), .ZN(n76));
  XNOR2_X1  g004(.A(69), .B(65), .ZN(n77));
  XNOR2_X1  g005(.A(77), .B(73), .ZN(n78));
  XNOR2_X1  g006(.A(n78), .B(n77), .ZN(n79));
  XNOR2_X1  g007(.A(85), .B(81), .ZN(n80));
  XNOR2_X1  g008(.A(93), .B(89), .ZN(n81));
  XNOR2_X1  g009(.A(n81), .B(n80), .ZN(n82));
  XNOR2_X1  g010(.A(n82), .B(n79), .ZN(n83));
  XNOR2_X1  g011(.A(n83), .B(n76), .ZN(n84));
  XNOR2_X1  g012(.A(n84), .B(n75), .ZN(n85));
  XOR2_X1   g013(.A(n84), .B(n75), .Z(n86));
  XNOR2_X1  g014(.A(29), .B(13), .ZN(n87));
  XNOR2_X1  g015(.A(61), .B(45), .ZN(n88));
  XNOR2_X1  g016(.A(n88), .B(n87), .ZN(n89));
  NAND2_X1  g017(.A1(137), .A2(132), .ZN(n90));
  XNOR2_X1  g018(.A(117), .B(113), .ZN(n91));
  XNOR2_X1  g019(.A(125), .B(121), .ZN(n92));
  XNOR2_X1  g020(.A(n92), .B(n91), .ZN(n93));
  XNOR2_X1  g021(.A(n93), .B(n82), .ZN(n94));
  XNOR2_X1  g022(.A(n94), .B(n90), .ZN(n95));
  XOR2_X1   g023(.A(n95), .B(n89), .Z(n96));
  XNOR2_X1  g024(.A(25), .B(9), .ZN(n97));
  XNOR2_X1  g025(.A(57), .B(41), .ZN(n98));
  XNOR2_X1  g026(.A(n98), .B(n97), .ZN(n99));
  NAND2_X1  g027(.A1(137), .A2(131), .ZN(n100));
  XNOR2_X1  g028(.A(101), .B(97), .ZN(n101));
  XNOR2_X1  g029(.A(109), .B(105), .ZN(n102));
  XNOR2_X1  g030(.A(n102), .B(n101), .ZN(n103));
  XNOR2_X1  g031(.A(n103), .B(n79), .ZN(n104));
  XNOR2_X1  g032(.A(n104), .B(n100), .ZN(n105));
  XOR2_X1   g033(.A(n105), .B(n99), .Z(n106));
  XNOR2_X1  g034(.A(21), .B(5), .ZN(n107));
  XNOR2_X1  g035(.A(53), .B(37), .ZN(n108));
  XNOR2_X1  g036(.A(n108), .B(n107), .ZN(n109));
  NAND2_X1  g037(.A1(137), .A2(130), .ZN(n110));
  XNOR2_X1  g038(.A(n103), .B(n93), .ZN(n111));
  XNOR2_X1  g039(.A(n111), .B(n110), .ZN(n112));
  XNOR2_X1  g040(.A(n112), .B(n109), .ZN(n113));
  NOR4_X1   g041(.A1(n106), .A2(n96), .A3(n86), .A4(n113), .ZN(n114));
  XOR2_X1   g042(.A(n112), .B(n109), .Z(n115));
  NOR4_X1   g043(.A1(n106), .A2(n96), .A3(n85), .A4(n115), .ZN(n116));
  XNOR2_X1  g044(.A(n95), .B(n89), .ZN(n117));
  NOR4_X1   g045(.A1(n106), .A2(n117), .A3(n86), .A4(n115), .ZN(n118));
  XNOR2_X1  g046(.A(n105), .B(n99), .ZN(n119));
  NOR4_X1   g047(.A1(n119), .A2(n96), .A3(n86), .A4(n115), .ZN(n120));
  NOR4_X1   g048(.A1(n118), .A2(n116), .A3(n114), .A4(n120), .ZN(n121));
  XNOR2_X1  g049(.A(81), .B(65), .ZN(n122));
  XNOR2_X1  g050(.A(113), .B(97), .ZN(n123));
  XNOR2_X1  g051(.A(n123), .B(n122), .ZN(n124));
  NAND2_X1  g052(.A1(137), .A2(133), .ZN(n125));
  XNOR2_X1  g053(.A(21), .B(17), .ZN(n126));
  XNOR2_X1  g054(.A(29), .B(25), .ZN(n127));
  XNOR2_X1  g055(.A(n127), .B(n126), .ZN(n128));
  XNOR2_X1  g056(.A(5), .B(\1 ), .ZN(n129));
  XNOR2_X1  g057(.A(13), .B(9), .ZN(n130));
  XNOR2_X1  g058(.A(n130), .B(n129), .ZN(n131));
  XNOR2_X1  g059(.A(n131), .B(n128), .ZN(n132));
  XNOR2_X1  g060(.A(n132), .B(n125), .ZN(n133));
  XOR2_X1   g061(.A(n133), .B(n124), .Z(n134));
  XNOR2_X1  g062(.A(85), .B(69), .ZN(n135));
  XNOR2_X1  g063(.A(117), .B(101), .ZN(n136));
  XNOR2_X1  g064(.A(n136), .B(n135), .ZN(n137));
  NAND2_X1  g065(.A1(137), .A2(134), .ZN(n138));
  XNOR2_X1  g066(.A(53), .B(49), .ZN(n139));
  XNOR2_X1  g067(.A(61), .B(57), .ZN(n140));
  XNOR2_X1  g068(.A(n140), .B(n139), .ZN(n141));
  XNOR2_X1  g069(.A(37), .B(33), .ZN(n142));
  XNOR2_X1  g070(.A(45), .B(41), .ZN(n143));
  XNOR2_X1  g071(.A(n143), .B(n142), .ZN(n144));
  XNOR2_X1  g072(.A(n144), .B(n141), .ZN(n145));
  XNOR2_X1  g073(.A(n145), .B(n138), .ZN(n146));
  XNOR2_X1  g074(.A(n146), .B(n137), .ZN(n147));
  NAND2_X1  g075(.A1(n147), .A2(n134), .ZN(n148));
  XNOR2_X1  g076(.A(93), .B(77), .ZN(n149));
  XNOR2_X1  g077(.A(125), .B(109), .ZN(n150));
  XNOR2_X1  g078(.A(n150), .B(n149), .ZN(n151));
  NAND2_X1  g079(.A1(137), .A2(136), .ZN(n152));
  XNOR2_X1  g080(.A(n141), .B(n128), .ZN(n153));
  XNOR2_X1  g081(.A(n153), .B(n152), .ZN(n154));
  XNOR2_X1  g082(.A(n154), .B(n151), .ZN(n155));
  XNOR2_X1  g083(.A(89), .B(73), .ZN(n156));
  XNOR2_X1  g084(.A(121), .B(105), .ZN(n157));
  XNOR2_X1  g085(.A(n157), .B(n156), .ZN(n158));
  NAND2_X1  g086(.A1(137), .A2(135), .ZN(n159));
  XNOR2_X1  g087(.A(n144), .B(n131), .ZN(n160));
  XNOR2_X1  g088(.A(n160), .B(n159), .ZN(n161));
  XOR2_X1   g089(.A(n161), .B(n158), .Z(n162));
  NAND2_X1  g090(.A1(n162), .A2(n155), .ZN(n163));
  OR4_X1    g091(.A1(n148), .A2(n121), .A3(n85), .A4(n163), .ZN(n164));
  XNOR2_X1  g092(.A(n164), .B(\1 ), .ZN(724));
  OR4_X1    g093(.A1(n148), .A2(n121), .A3(n113), .A4(n163), .ZN(n166));
  XNOR2_X1  g094(.A(n166), .B(5), .ZN(725));
  OR4_X1    g095(.A1(n148), .A2(n121), .A3(n119), .A4(n163), .ZN(n168));
  XNOR2_X1  g096(.A(n168), .B(9), .ZN(726));
  OR4_X1    g097(.A1(n148), .A2(n121), .A3(n117), .A4(n163), .ZN(n170));
  XNOR2_X1  g098(.A(n170), .B(13), .ZN(727));
  XNOR2_X1  g099(.A(n161), .B(n158), .ZN(n172));
  NAND3_X1  g100(.A1(n172), .A2(n147), .A3(n134), .ZN(n173));
  OR4_X1    g101(.A1(n155), .A2(n121), .A3(n85), .A4(n173), .ZN(n174));
  XNOR2_X1  g102(.A(n174), .B(17), .ZN(728));
  OR4_X1    g103(.A1(n155), .A2(n121), .A3(n113), .A4(n173), .ZN(n176));
  XNOR2_X1  g104(.A(n176), .B(21), .ZN(729));
  OR4_X1    g105(.A1(n155), .A2(n121), .A3(n119), .A4(n173), .ZN(n178));
  XNOR2_X1  g106(.A(n178), .B(25), .ZN(730));
  OR4_X1    g107(.A1(n155), .A2(n121), .A3(n117), .A4(n173), .ZN(n180));
  XNOR2_X1  g108(.A(n180), .B(29), .ZN(731));
  XNOR2_X1  g109(.A(n133), .B(n124), .ZN(n182));
  XOR2_X1   g110(.A(n146), .B(n137), .Z(n183));
  NAND2_X1  g111(.A1(n183), .A2(n182), .ZN(n184));
  OR4_X1    g112(.A1(n163), .A2(n121), .A3(n85), .A4(n184), .ZN(n185));
  XNOR2_X1  g113(.A(n185), .B(33), .ZN(732));
  OR4_X1    g114(.A1(n163), .A2(n121), .A3(n113), .A4(n184), .ZN(n187));
  XNOR2_X1  g115(.A(n187), .B(37), .ZN(733));
  OR4_X1    g116(.A1(n163), .A2(n121), .A3(n119), .A4(n184), .ZN(n189));
  XNOR2_X1  g117(.A(n189), .B(41), .ZN(734));
  OR4_X1    g118(.A1(n163), .A2(n121), .A3(n117), .A4(n184), .ZN(n191));
  XNOR2_X1  g119(.A(n191), .B(45), .ZN(735));
  NAND3_X1  g120(.A1(n172), .A2(n183), .A3(n182), .ZN(n193));
  OR4_X1    g121(.A1(n155), .A2(n121), .A3(n85), .A4(n193), .ZN(n194));
  XNOR2_X1  g122(.A(n194), .B(49), .ZN(736));
  OR4_X1    g123(.A1(n155), .A2(n121), .A3(n113), .A4(n193), .ZN(n196));
  XNOR2_X1  g124(.A(n196), .B(53), .ZN(737));
  OR4_X1    g125(.A1(n155), .A2(n121), .A3(n119), .A4(n193), .ZN(n198));
  XNOR2_X1  g126(.A(n198), .B(57), .ZN(738));
  OR4_X1    g127(.A1(n155), .A2(n121), .A3(n117), .A4(n193), .ZN(n200));
  XNOR2_X1  g128(.A(n200), .B(61), .ZN(739));
  NAND2_X1  g129(.A1(n113), .A2(n86), .ZN(n202));
  NAND2_X1  g130(.A1(n106), .A2(n117), .ZN(n203));
  XOR2_X1   g131(.A(n154), .B(n151), .Z(n204));
  NOR4_X1   g132(.A1(n204), .A2(n147), .A3(n134), .A4(n162), .ZN(n205));
  NOR4_X1   g133(.A1(n204), .A2(n183), .A3(n182), .A4(n162), .ZN(n206));
  NOR4_X1   g134(.A1(n155), .A2(n183), .A3(n134), .A4(n162), .ZN(n207));
  NOR4_X1   g135(.A1(n204), .A2(n183), .A3(n134), .A4(n172), .ZN(n208));
  NOR4_X1   g136(.A1(n207), .A2(n206), .A3(n205), .A4(n208), .ZN(n209));
  OR4_X1    g137(.A1(n182), .A2(n203), .A3(n202), .A4(n209), .ZN(n210));
  XNOR2_X1  g138(.A(n210), .B(65), .ZN(740));
  OR4_X1    g139(.A1(n147), .A2(n203), .A3(n202), .A4(n209), .ZN(n212));
  XNOR2_X1  g140(.A(n212), .B(69), .ZN(741));
  OR4_X1    g141(.A1(n172), .A2(n203), .A3(n202), .A4(n209), .ZN(n214));
  XNOR2_X1  g142(.A(n214), .B(73), .ZN(742));
  OR4_X1    g143(.A1(n155), .A2(n203), .A3(n202), .A4(n209), .ZN(n216));
  XNOR2_X1  g144(.A(n216), .B(77), .ZN(743));
  NAND3_X1  g145(.A1(n113), .A2(n119), .A3(n86), .ZN(n218));
  OR4_X1    g146(.A1(n182), .A2(n218), .A3(n117), .A4(n209), .ZN(n219));
  XNOR2_X1  g147(.A(n219), .B(81), .ZN(744));
  OR4_X1    g148(.A1(n147), .A2(n218), .A3(n117), .A4(n209), .ZN(n221));
  XNOR2_X1  g149(.A(n221), .B(85), .ZN(745));
  OR4_X1    g150(.A1(n172), .A2(n218), .A3(n117), .A4(n209), .ZN(n223));
  XNOR2_X1  g151(.A(n223), .B(89), .ZN(746));
  OR4_X1    g152(.A1(n155), .A2(n218), .A3(n117), .A4(n209), .ZN(n225));
  XNOR2_X1  g153(.A(n225), .B(93), .ZN(747));
  NAND2_X1  g154(.A1(n115), .A2(n85), .ZN(n227));
  OR4_X1    g155(.A1(n182), .A2(n203), .A3(n227), .A4(n209), .ZN(n228));
  XNOR2_X1  g156(.A(n228), .B(97), .ZN(748));
  OR4_X1    g157(.A1(n147), .A2(n203), .A3(n227), .A4(n209), .ZN(n230));
  XNOR2_X1  g158(.A(n230), .B(101), .ZN(749));
  OR4_X1    g159(.A1(n172), .A2(n203), .A3(n227), .A4(n209), .ZN(n232));
  XNOR2_X1  g160(.A(n232), .B(105), .ZN(750));
  OR4_X1    g161(.A1(n155), .A2(n203), .A3(n227), .A4(n209), .ZN(n234));
  XNOR2_X1  g162(.A(n234), .B(109), .ZN(751));
  NAND3_X1  g163(.A1(n115), .A2(n119), .A3(n85), .ZN(n236));
  OR4_X1    g164(.A1(n182), .A2(n236), .A3(n117), .A4(n209), .ZN(n237));
  XNOR2_X1  g165(.A(n237), .B(113), .ZN(752));
  OR4_X1    g166(.A1(n147), .A2(n236), .A3(n117), .A4(n209), .ZN(n239));
  XNOR2_X1  g167(.A(n239), .B(117), .ZN(753));
  OR4_X1    g168(.A1(n172), .A2(n236), .A3(n117), .A4(n209), .ZN(n241));
  XNOR2_X1  g169(.A(n241), .B(121), .ZN(754));
  OR4_X1    g170(.A1(n155), .A2(n236), .A3(n117), .A4(n209), .ZN(n243));
  XNOR2_X1  g171(.A(n243), .B(125), .ZN(755));
endmodule


