// Benchmark "c5315" written by ABC on Wed Oct 05 14:33:01 2022

module c5315 ( 
    \1 , 4, 11, 14, 17, 20, 23, 24, 25, 26, 27, 31, 34, 37, 40, 43, 46, 49,
    52, 53, 54, 61, 64, 67, 70, 73, 76, 79, 80, 81, 82, 83, 86, 87, 88, 91,
    94, 97, 100, 103, 106, 109, 112, 113, 114, 115, 116, 117, 118, 119,
    120, 121, 122, 123, 126, 127, 128, 129, 130, 131, 132, 135, 136, 137,
    140, 141, 145, 146, 149, 152, 155, 158, 161, 164, 167, 170, 173, 176,
    179, 182, 185, 188, 191, 194, 197, 200, 203, 206, 209, 210, 217, 218,
    225, 226, 233, 234, 241, 242, 245, 248, 251, 254, 257, 264, 265, 272,
    273, 280, 281, 288, 289, 292, 293, 299, 302, 307, 308, 315, 316, 323,
    324, 331, 332, 335, 338, 341, 348, 351, 358, 361, 366, 369, 372, 373,
    374, 386, 389, 400, 411, 422, 435, 446, 457, 468, 479, 490, 503, 514,
    523, 534, 545, 549, 552, 556, 559, 562, 566, 571, 574, 577, 580, 583,
    588, 591, 592, 595, 596, 597, 598, 599, 603, 607, 610, 613, 616, 619,
    625, 631,
    709, 816, 1066, 1137, 1138, 1139, 1140, 1141, 1142, 1143, 1144, 1145,
    1147, 1152, 1153, 1154, 1155, 1972, 2054, 2060, 2061, 2139, 2142, 2309,
    2387, 2527, 2584, 2590, 2623, 3357, 3358, 3359, 3360, 3604, 3613, 4272,
    4275, 4278, 4279, 4737, 4738, 4739, 4740, 5240, 5388, 6641, 6643, 6646,
    6648, 6716, 6877, 6924, 6925, 6926, 6927, 7015, 7363, 7365, 7432, 7449,
    7465, 7466, 7467, 7469, 7470, 7471, 7472, 7473, 7474, 7476, 7503, 7504,
    7506, 7511, 7515, 7516, 7517, 7518, 7519, 7520, 7521, 7522, 7600, 7601,
    7602, 7603, 7604, 7605, 7606, 7607, 7626, 7698, 7699, 7700, 7701, 7702,
    7703, 7704, 7705, 7706, 7707, 7735, 7736, 7737, 7738, 7739, 7740, 7741,
    7742, 7754, 7755, 7756, 7757, 7758, 7759, 7760, 7761, 8075, 8076, 8123,
    8124, 8127, 8128  );
  input  \1 , 4, 11, 14, 17, 20, 23, 24, 25, 26, 27, 31, 34, 37, 40, 43,
    46, 49, 52, 53, 54, 61, 64, 67, 70, 73, 76, 79, 80, 81, 82, 83, 86, 87,
    88, 91, 94, 97, 100, 103, 106, 109, 112, 113, 114, 115, 116, 117, 118,
    119, 120, 121, 122, 123, 126, 127, 128, 129, 130, 131, 132, 135, 136,
    137, 140, 141, 145, 146, 149, 152, 155, 158, 161, 164, 167, 170, 173,
    176, 179, 182, 185, 188, 191, 194, 197, 200, 203, 206, 209, 210, 217,
    218, 225, 226, 233, 234, 241, 242, 245, 248, 251, 254, 257, 264, 265,
    272, 273, 280, 281, 288, 289, 292, 293, 299, 302, 307, 308, 315, 316,
    323, 324, 331, 332, 335, 338, 341, 348, 351, 358, 361, 366, 369, 372,
    373, 374, 386, 389, 400, 411, 422, 435, 446, 457, 468, 479, 490, 503,
    514, 523, 534, 545, 549, 552, 556, 559, 562, 566, 571, 574, 577, 580,
    583, 588, 591, 592, 595, 596, 597, 598, 599, 603, 607, 610, 613, 616,
    619, 625, 631;
  output 709, 816, 1066, 1137, 1138, 1139, 1140, 1141, 1142, 1143, 1144, 1145,
    1147, 1152, 1153, 1154, 1155, 1972, 2054, 2060, 2061, 2139, 2142, 2309,
    2387, 2527, 2584, 2590, 2623, 3357, 3358, 3359, 3360, 3604, 3613, 4272,
    4275, 4278, 4279, 4737, 4738, 4739, 4740, 5240, 5388, 6641, 6643, 6646,
    6648, 6716, 6877, 6924, 6925, 6926, 6927, 7015, 7363, 7365, 7432, 7449,
    7465, 7466, 7467, 7469, 7470, 7471, 7472, 7473, 7474, 7476, 7503, 7504,
    7506, 7511, 7515, 7516, 7517, 7518, 7519, 7520, 7521, 7522, 7600, 7601,
    7602, 7603, 7604, 7605, 7606, 7607, 7626, 7698, 7699, 7700, 7701, 7702,
    7703, 7704, 7705, 7706, 7707, 7735, 7736, 7737, 7738, 7739, 7740, 7741,
    7742, 7754, 7755, 7756, 7757, 7758, 7759, 7760, 7761, 8075, 8076, 8123,
    8124, 8127, 8128;
  wire n314, n316, n322, n324, n327, n328, n329, n330, n332, n333, n335,
    n336, n338, n339, n341, n342, n343, n344, n345, n346, n347, n348, n349,
    n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
    n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
    n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
    n386, n387, n388, n390, n391, n392, n393, n394, n395, n396, n397, n398,
    n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
    n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
    n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
    n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
    n447, n448, n449, n450, n451, n452, n453, n455, n456, n457, n458, n459,
    n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
    n472, n473, n474, n475, n476, n477, n479, n480, n481, n482, n483, n484,
    n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
    n497, n498, n499, n500, n502, n503, n506, n507, n508, n509, n510, n511,
    n512, n513, n514, n515, n516, n518, n519, n520, n521, n522, n523, n524,
    n525, n526, n527, n528, n529, n530, n531, n532, n534, n535, n536, n537,
    n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
    n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n561, n562,
    n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
    n575, n576, n577, n583, n584, n585, n586, n587, n588, n590, n591, n592,
    n593, n594, n595, n597, n598, n599, n600, n602, n603, n604, n605, n606,
    n607, n608, n609, n610, n612, n613, n614, n615, n616, n617, n619, n620,
    n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n632, n633,
    n634, n635, n637, n638, n639, n640, n641, n642, n644, n645, n646, n647,
    n648, n649, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
    n661, n663, n664, n665, n666, n667, n669, n670, n671, n672, n673, n674,
    n676, n677, n678, n679, n681, n682, n683, n684, n685, n686, n687, n688,
    n689, n690, n691, n692, n693, n694, n696, n697, n698, n699, n700, n701,
    n702, n703, n704, n705, n706, n707, n708, n709, n710, n712, n713, n714,
    n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
    n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n738, n739,
    n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
    n752, n754, n755, n756, n757, n758, n759, n760, n761, n762, n764, n765,
    n766, n767, n768, n769, n770, n771, n772, n774, n776, n778, n780, n782,
    n784, n786, n788, n790, n791, n793, n794, n796, n797, n799, n800, n802,
    n803, n804, n805, n807, n808, n809, n810, n812, n813, n814, n815, n817,
    n818, n819, n820, n822, n823, n824, n825, n826, n827, n828, n829, n830,
    n833, n834, n836, n837, n839, n840, n842, n843, n845, n846, n848, n850,
    n851, n853, n854, n856, n857, n859, n861, n863, n865, n867, n869, n871,
    n873, n875, n876, n878, n879, n881, n882, n884, n885, n887, n888, n889,
    n890, n892, n893, n894, n895, n897, n898, n899, n900, n902, n903, n904,
    n905, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
    n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
    n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n942,
    n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
    n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
    n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
    n979, n980, n981, n982, n983, n985, n986, n987, n988, n989, n990, n991,
    n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
    n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
    n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
    n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
    n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
    n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
    n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
    n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
    n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
    n1083, n1084, n1085, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
    n1095, n1097, n1098, n1100, n1101, n1102, n1103;
  INV_X1    g000(.A(545), .ZN(1137));
  INV_X1    g001(.A(348), .ZN(1138));
  INV_X1    g002(.A(366), .ZN(1139));
  AND2_X1   g003(.A1(562), .A2(552), .ZN(1140));
  INV_X1    g004(.A(549), .ZN(1141));
  INV_X1    g005(.A(338), .ZN(1144));
  INV_X1    g006(.A(358), .ZN(1145));
  AND2_X1   g007(.A1(145), .A2(141), .ZN(1147));
  INV_X1    g008(.A(245), .ZN(1152));
  INV_X1    g009(.A(552), .ZN(1153));
  INV_X1    g010(.A(562), .ZN(1154));
  INV_X1    g011(.A(559), .ZN(1155));
  AND2_X1   g012(.A1(373), .A2(\1 ), .ZN(1972));
  INV_X1    g013(.A(136), .ZN(n314));
  NOR2_X1   g014(.A1(592), .A2(n314), .ZN(2054));
  INV_X1    g015(.A(591), .ZN(n316));
  NAND2_X1  g016(.A1(n316), .A2(27), .ZN(2060));
  NAND2_X1  g017(.A1(556), .A2(386), .ZN(2061));
  NAND3_X1  g018(.A1(140), .A2(31), .A3(27), .ZN(2590));
  NAND2_X1  g019(.A1(31), .A2(27), .ZN(2623));
  INV_X1    g020(.A(299), .ZN(3613));
  MUX2_X1   g021(.S(588), .B(87), .A(86), .ZN(n322));
  NAND3_X1  g022(.A1(n322), .A2(31), .A3(27), .ZN(4272));
  MUX2_X1   g023(.S(588), .B(34), .A(88), .ZN(n324));
  NAND3_X1  g024(.A1(n324), .A2(31), .A3(27), .ZN(4275));
  NAND3_X1  g025(.A1(83), .A2(31), .A3(27), .ZN(4279));
  INV_X1    g026(.A(141), .ZN(n327));
  INV_X1    g027(.A(588), .ZN(n328));
  AND4_X1   g028(.A1(31), .A2(27), .A3(25), .A4(588), .ZN(n329));
  AOI211_X1 g029(.A(2623), .B(n329), .C1(n328), .C2(24), .ZN(n330));
  NOR2_X1   g030(.A1(n330), .A2(n327), .ZN(4737));
  AND4_X1   g031(.A1(81), .A2(31), .A3(27), .A4(588), .ZN(n332));
  AOI211_X1 g032(.A(2623), .B(n332), .C1(n328), .C2(26), .ZN(n333));
  NOR2_X1   g033(.A1(n333), .A2(n327), .ZN(4738));
  AND4_X1   g034(.A1(31), .A2(27), .A3(23), .A4(588), .ZN(n335));
  AOI211_X1 g035(.A(2623), .B(n335), .C1(n328), .C2(79), .ZN(n336));
  NOR2_X1   g036(.A1(n336), .A2(n327), .ZN(4739));
  AND4_X1   g037(.A1(80), .A2(31), .A3(27), .A4(588), .ZN(n338));
  AOI211_X1 g038(.A(2623), .B(n338), .C1(n328), .C2(82), .ZN(n339));
  NOR2_X1   g039(.A1(n339), .A2(n327), .ZN(4740));
  INV_X1    g040(.A(595), .ZN(n341));
  NOR2_X1   g041(.A1(596), .A2(341), .ZN(n342));
  AOI211_X1 g042(.A(523), .B(n342), .C1(n341), .C2(341), .ZN(n343));
  INV_X1    g043(.A(341), .ZN(n344));
  INV_X1    g044(.A(523), .ZN(n345));
  NOR3_X1   g045(.A1(598), .A2(n345), .A3(n344), .ZN(n346));
  NOR3_X1   g046(.A1(597), .A2(n345), .A3(341), .ZN(n347));
  NOR3_X1   g047(.A1(n347), .A2(n346), .A3(n343), .ZN(n348));
  INV_X1    g048(.A(248), .ZN(n349));
  INV_X1    g049(.A(251), .ZN(n350));
  INV_X1    g050(.A(361), .ZN(n351));
  MUX2_X1   g051(.S(n351), .B(n350), .A(n349), .ZN(n352));
  INV_X1    g052(.A(302), .ZN(n353));
  MUX2_X1   g053(.S(n353), .B(n350), .A(n349), .ZN(n354));
  INV_X1    g054(.A(242), .ZN(n355));
  INV_X1    g055(.A(254), .ZN(n356));
  INV_X1    g056(.A(293), .ZN(n357));
  MUX2_X1   g057(.S(n357), .B(n356), .A(n355), .ZN(n358));
  INV_X1    g058(.A(n358), .ZN(n359));
  MUX2_X1   g059(.S(514), .B(598), .A(n341), .ZN(n360));
  OR4_X1    g060(.A1(n359), .A2(n354), .A3(n352), .A4(n360), .ZN(n361));
  INV_X1    g061(.A(490), .ZN(n362));
  OAI21_X1  g062(.A(n362), .B1(316), .B2(n356), .ZN(n363));
  AOI21_X1  g063(.A(n363), .B1(316), .B2(242), .ZN(n364));
  AND3_X1   g064(.A1(490), .A2(316), .A3(248), .ZN(n365));
  NOR3_X1   g065(.A1(n362), .A2(316), .A3(n350), .ZN(n366));
  NOR3_X1   g066(.A1(n366), .A2(n365), .A3(n364), .ZN(n367));
  NOR2_X1   g067(.A1(596), .A2(324), .ZN(n368));
  AOI211_X1 g068(.A(503), .B(n368), .C1(n341), .C2(324), .ZN(n369));
  INV_X1    g069(.A(324), .ZN(n370));
  INV_X1    g070(.A(503), .ZN(n371));
  NOR3_X1   g071(.A1(598), .A2(n371), .A3(n370), .ZN(n372));
  NOR3_X1   g072(.A1(597), .A2(n371), .A3(324), .ZN(n373));
  NOR3_X1   g073(.A1(n373), .A2(n372), .A3(n369), .ZN(n374));
  INV_X1    g074(.A(479), .ZN(n375));
  OAI21_X1  g075(.A(n375), .B1(308), .B2(n356), .ZN(n376));
  AOI21_X1  g076(.A(n376), .B1(308), .B2(242), .ZN(n377));
  AND3_X1   g077(.A1(479), .A2(308), .A3(248), .ZN(n378));
  NOR3_X1   g078(.A1(n375), .A2(308), .A3(n350), .ZN(n379));
  NOR3_X1   g079(.A1(n379), .A2(n378), .A3(n377), .ZN(n380));
  NOR2_X1   g080(.A1(596), .A2(351), .ZN(n381));
  AOI211_X1 g081(.A(534), .B(n381), .C1(n341), .C2(351), .ZN(n382));
  INV_X1    g082(.A(351), .ZN(n383));
  INV_X1    g083(.A(534), .ZN(n384));
  NOR3_X1   g084(.A1(598), .A2(n384), .A3(n383), .ZN(n385));
  NOR3_X1   g085(.A1(597), .A2(n384), .A3(351), .ZN(n386));
  NOR3_X1   g086(.A1(n386), .A2(n385), .A3(n382), .ZN(n387));
  OR4_X1    g087(.A1(n380), .A2(n374), .A3(n367), .A4(n387), .ZN(n388));
  NOR3_X1   g088(.A1(n388), .A2(n361), .A3(n348), .ZN(5240));
  INV_X1    g089(.A(446), .ZN(n390));
  OAI21_X1  g090(.A(n390), .B1(n356), .B2(206), .ZN(n391));
  AOI21_X1  g091(.A(n391), .B1(242), .B2(206), .ZN(n392));
  AND3_X1   g092(.A1(446), .A2(248), .A3(206), .ZN(n393));
  NOR3_X1   g093(.A1(n390), .A2(n350), .A3(206), .ZN(n394));
  NOR3_X1   g094(.A1(n394), .A2(n393), .A3(n392), .ZN(n395));
  NOR2_X1   g095(.A1(596), .A2(210), .ZN(n396));
  AOI211_X1 g096(.A(457), .B(n396), .C1(n341), .C2(210), .ZN(n397));
  INV_X1    g097(.A(210), .ZN(n398));
  INV_X1    g098(.A(457), .ZN(n399));
  NOR3_X1   g099(.A1(598), .A2(n399), .A3(n398), .ZN(n400));
  NOR3_X1   g100(.A1(597), .A2(n399), .A3(210), .ZN(n401));
  NOR3_X1   g101(.A1(n401), .A2(n400), .A3(n397), .ZN(n402));
  NOR2_X1   g102(.A1(596), .A2(218), .ZN(n403));
  AOI211_X1 g103(.A(468), .B(n403), .C1(n341), .C2(218), .ZN(n404));
  INV_X1    g104(.A(218), .ZN(n405));
  INV_X1    g105(.A(468), .ZN(n406));
  NOR3_X1   g106(.A1(598), .A2(n406), .A3(n405), .ZN(n407));
  NOR3_X1   g107(.A1(597), .A2(n406), .A3(218), .ZN(n408));
  NOR3_X1   g108(.A1(n408), .A2(n407), .A3(n404), .ZN(n409));
  OR3_X1    g109(.A1(n409), .A2(n402), .A3(n395), .ZN(n410));
  NOR2_X1   g110(.A1(596), .A2(281), .ZN(n411));
  AOI211_X1 g111(.A(374), .B(n411), .C1(n341), .C2(281), .ZN(n412));
  INV_X1    g112(.A(281), .ZN(n413));
  INV_X1    g113(.A(374), .ZN(n414));
  NOR3_X1   g114(.A1(598), .A2(n414), .A3(n413), .ZN(n415));
  NOR3_X1   g115(.A1(597), .A2(n414), .A3(281), .ZN(n416));
  NOR3_X1   g116(.A1(n416), .A2(n415), .A3(n412), .ZN(n417));
  NOR2_X1   g117(.A1(596), .A2(273), .ZN(n418));
  AOI211_X1 g118(.A(411), .B(n418), .C1(n341), .C2(273), .ZN(n419));
  INV_X1    g119(.A(273), .ZN(n420));
  INV_X1    g120(.A(411), .ZN(n421));
  NOR3_X1   g121(.A1(598), .A2(n421), .A3(n420), .ZN(n422));
  NOR3_X1   g122(.A1(597), .A2(n421), .A3(273), .ZN(n423));
  NOR3_X1   g123(.A1(n423), .A2(n422), .A3(n419), .ZN(n424));
  NOR2_X1   g124(.A1(596), .A2(257), .ZN(n425));
  AOI211_X1 g125(.A(389), .B(n425), .C1(n341), .C2(257), .ZN(n426));
  INV_X1    g126(.A(257), .ZN(n427));
  INV_X1    g127(.A(389), .ZN(n428));
  NOR3_X1   g128(.A1(598), .A2(n428), .A3(n427), .ZN(n429));
  NOR3_X1   g129(.A1(597), .A2(n428), .A3(257), .ZN(n430));
  NOR3_X1   g130(.A1(n430), .A2(n429), .A3(n426), .ZN(n431));
  NOR2_X1   g131(.A1(596), .A2(265), .ZN(n432));
  AOI211_X1 g132(.A(400), .B(n432), .C1(n341), .C2(265), .ZN(n433));
  INV_X1    g133(.A(265), .ZN(n434));
  INV_X1    g134(.A(400), .ZN(n435));
  NOR3_X1   g135(.A1(598), .A2(n435), .A3(n434), .ZN(n436));
  NOR3_X1   g136(.A1(597), .A2(n435), .A3(265), .ZN(n437));
  NOR3_X1   g137(.A1(n437), .A2(n436), .A3(n433), .ZN(n438));
  NOR2_X1   g138(.A1(596), .A2(234), .ZN(n439));
  AOI211_X1 g139(.A(435), .B(n439), .C1(n341), .C2(234), .ZN(n440));
  INV_X1    g140(.A(234), .ZN(n441));
  INV_X1    g141(.A(435), .ZN(n442));
  NOR3_X1   g142(.A1(598), .A2(n442), .A3(n441), .ZN(n443));
  NOR3_X1   g143(.A1(597), .A2(n442), .A3(234), .ZN(n444));
  NOR3_X1   g144(.A1(n444), .A2(n443), .A3(n440), .ZN(n445));
  NOR2_X1   g145(.A1(596), .A2(226), .ZN(n446));
  AOI211_X1 g146(.A(422), .B(n446), .C1(n341), .C2(226), .ZN(n447));
  INV_X1    g147(.A(226), .ZN(n448));
  INV_X1    g148(.A(422), .ZN(n449));
  NOR3_X1   g149(.A1(598), .A2(n449), .A3(n448), .ZN(n450));
  NOR3_X1   g150(.A1(597), .A2(n449), .A3(226), .ZN(n451));
  NOR3_X1   g151(.A1(n451), .A2(n450), .A3(n447), .ZN(n452));
  OR4_X1    g152(.A1(n445), .A2(n438), .A3(n431), .A4(n452), .ZN(n453));
  NOR4_X1   g153(.A1(n424), .A2(n417), .A3(n410), .A4(n453), .ZN(5388));
  MUX2_X1   g154(.S(335), .B(209), .A(206), .ZN(n455));
  XNOR2_X1  g155(.A(n455), .B(446), .ZN(n456));
  INV_X1    g156(.A(n456), .ZN(n457));
  MUX2_X1   g157(.S(335), .B(217), .A(210), .ZN(n458));
  XNOR2_X1  g158(.A(n458), .B(n399), .ZN(n459));
  MUX2_X1   g159(.S(335), .B(233), .A(226), .ZN(n460));
  XNOR2_X1  g160(.A(n460), .B(422), .ZN(n461));
  MUX2_X1   g161(.S(335), .B(225), .A(218), .ZN(n462));
  XNOR2_X1  g162(.A(n462), .B(468), .ZN(n463));
  NOR2_X1   g163(.A1(n463), .A2(n461), .ZN(n464));
  MUX2_X1   g164(.S(335), .B(288), .A(281), .ZN(n465));
  XNOR2_X1  g165(.A(n465), .B(374), .ZN(n466));
  MUX2_X1   g166(.S(335), .B(280), .A(273), .ZN(n467));
  XNOR2_X1  g167(.A(n467), .B(411), .ZN(n468));
  NOR2_X1   g168(.A1(n468), .A2(n466), .ZN(n469));
  MUX2_X1   g169(.S(335), .B(272), .A(265), .ZN(n470));
  XNOR2_X1  g170(.A(n470), .B(n435), .ZN(n471));
  MUX2_X1   g171(.S(335), .B(241), .A(234), .ZN(n472));
  XNOR2_X1  g172(.A(n472), .B(435), .ZN(n473));
  INV_X1    g173(.A(n473), .ZN(n474));
  MUX2_X1   g174(.S(335), .B(264), .A(257), .ZN(n475));
  XNOR2_X1  g175(.A(n475), .B(n428), .ZN(n476));
  AND4_X1   g176(.A1(n474), .A2(n471), .A3(n469), .A4(n476), .ZN(n477));
  AND4_X1   g177(.A1(n464), .A2(n459), .A3(n457), .A4(n477), .ZN(6641));
  MUX2_X1   g178(.S(332), .B(315), .A(308), .ZN(n479));
  XNOR2_X1  g179(.A(n479), .B(n375), .ZN(n480));
  MUX2_X1   g180(.S(332), .B(323), .A(316), .ZN(n481));
  XNOR2_X1  g181(.A(n481), .B(n362), .ZN(n482));
  MUX2_X1   g182(.S(332), .B(3613), .A(n357), .ZN(n483));
  INV_X1    g183(.A(307), .ZN(n484));
  MUX2_X1   g184(.S(332), .B(n484), .A(n353), .ZN(n485));
  NAND4_X1  g185(.A1(n483), .A2(n482), .A3(n480), .A4(n485), .ZN(n486));
  MUX2_X1   g186(.S(332), .B(358), .A(351), .ZN(n487));
  XNOR2_X1  g187(.A(n487), .B(534), .ZN(n488));
  MUX2_X1   g188(.S(332), .B(366), .A(361), .ZN(n489));
  NOR2_X1   g189(.A1(n489), .A2(n488), .ZN(n490));
  MUX2_X1   g190(.S(332), .B(331), .A(324), .ZN(n491));
  XNOR2_X1  g191(.A(n491), .B(503), .ZN(n492));
  INV_X1    g192(.A(n492), .ZN(n493));
  MUX2_X1   g193(.S(332), .B(348), .A(341), .ZN(n494));
  XNOR2_X1  g194(.A(n494), .B(523), .ZN(n495));
  INV_X1    g195(.A(n495), .ZN(n496));
  INV_X1    g196(.A(332), .ZN(n497));
  NOR2_X1   g197(.A1(338), .A2(n497), .ZN(n498));
  XNOR2_X1  g198(.A(n498), .B(514), .ZN(n499));
  NAND4_X1  g199(.A1(n496), .A2(n493), .A3(n490), .A4(n499), .ZN(n500));
  NOR2_X1   g200(.A1(n500), .A2(n486), .ZN(6643));
  AND3_X1   g201(.A1(n485), .A2(n482), .A3(n480), .ZN(n502));
  AND4_X1   g202(.A1(n496), .A2(n493), .A3(n490), .A4(n499), .ZN(n503));
  AND3_X1   g203(.A1(n503), .A2(n502), .A3(n483), .ZN(6646));
  AND4_X1   g204(.A1(n464), .A2(n459), .A3(n457), .A4(n477), .ZN(6648));
  XOR2_X1   g205(.A(316), .B(308), .ZN(n506));
  XNOR2_X1  g206(.A(302), .B(293), .ZN(n507));
  XNOR2_X1  g207(.A(n507), .B(n506), .ZN(n508));
  XNOR2_X1  g208(.A(369), .B(361), .ZN(n509));
  XNOR2_X1  g209(.A(351), .B(341), .ZN(n510));
  INV_X1    g210(.A(n510), .ZN(n511));
  NOR3_X1   g211(.A1(n511), .A2(n509), .A3(n370), .ZN(n512));
  NOR3_X1   g212(.A1(n510), .A2(n509), .A3(324), .ZN(n513));
  AND3_X1   g213(.A1(n510), .A2(n509), .A3(n370), .ZN(n514));
  AND3_X1   g214(.A1(n511), .A2(n509), .A3(324), .ZN(n515));
  NOR4_X1   g215(.A1(n514), .A2(n513), .A3(n512), .A4(n515), .ZN(n516));
  XNOR2_X1  g216(.A(n516), .B(n508), .ZN(6716));
  XNOR2_X1  g217(.A(226), .B(218), .ZN(n518));
  XNOR2_X1  g218(.A(210), .B(206), .ZN(n519));
  XNOR2_X1  g219(.A(n519), .B(n518), .ZN(n520));
  XNOR2_X1  g220(.A(289), .B(281), .ZN(n521));
  XNOR2_X1  g221(.A(257), .B(234), .ZN(n522));
  INV_X1    g222(.A(n522), .ZN(n523));
  XNOR2_X1  g223(.A(273), .B(265), .ZN(n524));
  INV_X1    g224(.A(n524), .ZN(n525));
  NOR3_X1   g225(.A1(n525), .A2(n523), .A3(n521), .ZN(n526));
  NOR3_X1   g226(.A1(n524), .A2(n522), .A3(n521), .ZN(n527));
  INV_X1    g227(.A(n521), .ZN(n528));
  NOR3_X1   g228(.A1(n525), .A2(n522), .A3(n528), .ZN(n529));
  NOR3_X1   g229(.A1(n524), .A2(n523), .A3(n528), .ZN(n530));
  NOR4_X1   g230(.A1(n529), .A2(n527), .A3(n526), .A4(n530), .ZN(n531));
  XNOR2_X1  g231(.A(n531), .B(n520), .ZN(n532));
  INV_X1    g232(.A(n532), .ZN(6877));
  NAND3_X1  g233(.A1(n464), .A2(n459), .A3(n457), .ZN(n534));
  INV_X1    g234(.A(n459), .ZN(n535));
  AND2_X1   g235(.A1(n462), .A2(468), .ZN(n536));
  INV_X1    g236(.A(n536), .ZN(n537));
  NOR3_X1   g237(.A1(n537), .A2(n535), .A3(n456), .ZN(n538));
  XNOR2_X1  g238(.A(n462), .B(n406), .ZN(n539));
  AND2_X1   g239(.A1(n460), .A2(422), .ZN(n540));
  AND4_X1   g240(.A1(n539), .A2(n459), .A3(n457), .A4(n540), .ZN(n541));
  AND2_X1   g241(.A1(n455), .A2(446), .ZN(n542));
  NAND2_X1  g242(.A1(n458), .A2(457), .ZN(n543));
  NOR2_X1   g243(.A1(n543), .A2(n456), .ZN(n544));
  NOR4_X1   g244(.A1(n542), .A2(n541), .A3(n538), .A4(n544), .ZN(n545));
  XNOR2_X1  g245(.A(n470), .B(400), .ZN(n546));
  NOR2_X1   g246(.A1(n546), .A2(n468), .ZN(n547));
  AND2_X1   g247(.A1(n465), .A2(374), .ZN(n548));
  AND4_X1   g248(.A1(n547), .A2(n476), .A3(n474), .A4(n548), .ZN(n549));
  XNOR2_X1  g249(.A(n475), .B(389), .ZN(n550));
  NAND2_X1  g250(.A1(n470), .A2(400), .ZN(n551));
  NOR3_X1   g251(.A1(n551), .A2(n550), .A3(n473), .ZN(n552));
  NAND2_X1  g252(.A1(n467), .A2(411), .ZN(n553));
  NOR4_X1   g253(.A1(n550), .A2(n473), .A3(n546), .A4(n553), .ZN(n554));
  AND2_X1   g254(.A1(n472), .A2(435), .ZN(n555));
  AND2_X1   g255(.A1(n475), .A2(389), .ZN(n556));
  AOI211_X1 g256(.A(n555), .B(n554), .C1(n474), .C2(n556), .ZN(n557));
  INV_X1    g257(.A(n557), .ZN(n558));
  NOR3_X1   g258(.A1(n558), .A2(n552), .A3(n549), .ZN(n559));
  OAI21_X1  g259(.A(n545), .B1(n559), .B2(n534), .ZN(6924));
  INV_X1    g260(.A(n483), .ZN(n561));
  INV_X1    g261(.A(n485), .ZN(n562));
  AND2_X1   g262(.A1(n481), .A2(490), .ZN(n563));
  AND4_X1   g263(.A1(n485), .A2(n483), .A3(n480), .A4(n563), .ZN(n564));
  AND2_X1   g264(.A1(n479), .A2(479), .ZN(n565));
  NOR4_X1   g265(.A1(n564), .A2(n562), .A3(n561), .A4(n565), .ZN(n566));
  NOR2_X1   g266(.A1(n495), .A2(n488), .ZN(n567));
  NAND4_X1  g267(.A1(n499), .A2(n493), .A3(n489), .A4(n567), .ZN(n568));
  AND2_X1   g268(.A1(n494), .A2(523), .ZN(n569));
  NAND3_X1  g269(.A1(n569), .A2(n499), .A3(n493), .ZN(n570));
  INV_X1    g270(.A(n499), .ZN(n571));
  NAND2_X1  g271(.A1(n487), .A2(534), .ZN(n572));
  OR4_X1    g272(.A1(n571), .A2(n495), .A3(n492), .A4(n572), .ZN(n573));
  OAI21_X1  g273(.A(514), .B1(338), .B2(n497), .ZN(n574));
  NOR2_X1   g274(.A1(n574), .A2(n492), .ZN(n575));
  AOI21_X1  g275(.A(n575), .B1(n491), .B2(503), .ZN(n576));
  AND4_X1   g276(.A1(n573), .A2(n570), .A3(n568), .A4(n576), .ZN(n577));
  OAI21_X1  g277(.A(n566), .B1(n577), .B2(n486), .ZN(6925));
  OAI21_X1  g278(.A(n545), .B1(n559), .B2(n534), .ZN(6926));
  OAI21_X1  g279(.A(n566), .B1(n577), .B2(n486), .ZN(6927));
  INV_X1    g280(.A(619), .ZN(n583));
  INV_X1    g281(.A(54), .ZN(n584));
  XNOR2_X1  g282(.A(n489), .B(n584), .ZN(n585));
  NOR3_X1   g283(.A1(n585), .A2(625), .A3(n583), .ZN(n586));
  AND3_X1   g284(.A1(625), .A2(n583), .A3(131), .ZN(n587));
  NOR2_X1   g285(.A1(625), .A2(619), .ZN(n588));
  AOI211_X1 g286(.A(n587), .B(n586), .C1(n352), .C2(n588), .ZN(7015));
  NOR2_X1   g287(.A1(625), .A2(n583), .ZN(n590));
  INV_X1    g288(.A(n590), .ZN(n591));
  NOR2_X1   g289(.A1(n489), .A2(54), .ZN(n592));
  XNOR2_X1  g290(.A(n592), .B(n488), .ZN(n593));
  NOR2_X1   g291(.A1(n593), .A2(n591), .ZN(n594));
  AND3_X1   g292(.A1(625), .A2(n583), .A3(129), .ZN(n595));
  AOI211_X1 g293(.A(n594), .B(n595), .C1(n588), .C2(n387), .ZN(7363));
  INV_X1    g294(.A(4), .ZN(n597));
  XNOR2_X1  g295(.A(n466), .B(n597), .ZN(n598));
  NOR2_X1   g296(.A1(n598), .A2(n591), .ZN(n599));
  AND3_X1   g297(.A1(625), .A2(n583), .A3(117), .ZN(n600));
  AOI211_X1 g298(.A(n599), .B(n600), .C1(n588), .C2(n417), .ZN(7365));
  OAI21_X1  g299(.A(n577), .B1(n500), .B2(n584), .ZN(n602));
  INV_X1    g300(.A(n565), .ZN(n603));
  NAND3_X1  g301(.A1(n563), .A2(n485), .A3(n480), .ZN(n604));
  NAND3_X1  g302(.A1(n604), .A2(n603), .A3(n485), .ZN(n605));
  XNOR2_X1  g303(.A(n605), .B(n561), .ZN(n606));
  INV_X1    g304(.A(n606), .ZN(n607));
  NAND2_X1  g305(.A1(n482), .A2(n480), .ZN(n608));
  AND4_X1   g306(.A1(n603), .A2(n608), .A3(n485), .A4(n604), .ZN(n609));
  XNOR2_X1  g307(.A(n609), .B(n561), .ZN(n610));
  MUX2_X1   g308(.S(n602), .B(n610), .A(n607), .ZN(7432));
  INV_X1    g309(.A(607), .ZN(n612));
  NAND2_X1  g310(.A1(610), .A2(n612), .ZN(n613));
  OR2_X1    g311(.A1(610), .A2(607), .ZN(n614));
  AND2_X1   g312(.A1(610), .A2(607), .ZN(n615));
  NOR2_X1   g313(.A1(610), .A2(n612), .ZN(n616));
  AOI22_X1  g314(.A1(n615), .A2(61), .B1(11), .B2(n616), .ZN(n617));
  OAI221_X1 g315(.A(n617), .B1(n613), .B2(7365), .C1(7015), .C2(n614), .ZN(7449));
  NOR4_X1   g316(.A1(n489), .A2(n488), .A3(n584), .A4(n495), .ZN(n619));
  MUX2_X1   g317(.S(332), .B(1139), .A(n351), .ZN(n620));
  NOR3_X1   g318(.A1(n495), .A2(n620), .A3(n488), .ZN(n621));
  NAND2_X1  g319(.A1(n621), .A2(n499), .ZN(n622));
  NOR2_X1   g320(.A1(n572), .A2(n495), .ZN(n623));
  NAND2_X1  g321(.A1(n623), .A2(n499), .ZN(n624));
  NAND2_X1  g322(.A1(n569), .A2(n499), .ZN(n625));
  NAND4_X1  g323(.A1(n624), .A2(n622), .A3(n574), .A4(n625), .ZN(n626));
  AOI21_X1  g324(.A(n626), .B1(n619), .B2(n499), .ZN(n627));
  XNOR2_X1  g325(.A(n627), .B(n492), .ZN(n628));
  INV_X1    g326(.A(n628), .ZN(n629));
  AND3_X1   g327(.A1(625), .A2(n583), .A3(52), .ZN(n630));
  AOI221_X1 g328(.A(n630), .B1(n588), .B2(n374), .C1(n590), .C2(n629), .ZN(7465));
  NOR4_X1   g329(.A1(n621), .A2(n619), .A3(n569), .A4(n623), .ZN(n632));
  XNOR2_X1  g330(.A(n632), .B(n571), .ZN(n633));
  NOR2_X1   g331(.A1(n633), .A2(n591), .ZN(n634));
  AND3_X1   g332(.A1(625), .A2(n583), .A3(130), .ZN(n635));
  AOI211_X1 g333(.A(n634), .B(n635), .C1(n588), .C2(n360), .ZN(7466));
  NOR3_X1   g334(.A1(n489), .A2(n488), .A3(n584), .ZN(n637));
  OAI21_X1  g335(.A(n572), .B1(n620), .B2(n488), .ZN(n638));
  NOR2_X1   g336(.A1(n638), .A2(n637), .ZN(n639));
  XNOR2_X1  g337(.A(n639), .B(n495), .ZN(n640));
  NOR2_X1   g338(.A1(n640), .A2(n591), .ZN(n641));
  AND3_X1   g339(.A1(625), .A2(n583), .A3(119), .ZN(n642));
  AOI211_X1 g340(.A(n641), .B(n642), .C1(n588), .C2(n348), .ZN(7467));
  INV_X1    g341(.A(616), .ZN(n644));
  NAND2_X1  g342(.A1(n644), .A2(613), .ZN(n645));
  OR2_X1    g343(.A1(616), .A2(613), .ZN(n646));
  AND2_X1   g344(.A1(616), .A2(613), .ZN(n647));
  NOR2_X1   g345(.A1(n644), .A2(613), .ZN(n648));
  AOI22_X1  g346(.A1(n647), .A2(61), .B1(11), .B2(n648), .ZN(n649));
  OAI221_X1 g347(.A(n649), .B1(n645), .B2(7365), .C1(7015), .C2(n646), .ZN(7469));
  NOR4_X1   g348(.A1(n468), .A2(n466), .A3(n597), .A4(n546), .ZN(n651));
  NAND2_X1  g349(.A1(n465), .A2(374), .ZN(n652));
  OR3_X1    g350(.A1(n652), .A2(n546), .A3(n468), .ZN(n653));
  OR3_X1    g351(.A1(n553), .A2(n550), .A3(n546), .ZN(n654));
  AND2_X1   g352(.A1(n470), .A2(400), .ZN(n655));
  AOI21_X1  g353(.A(n556), .B1(n655), .B2(n476), .ZN(n656));
  OAI211_X1 g354(.A(n654), .B(n656), .C1(n653), .C2(n550), .ZN(n657));
  AOI21_X1  g355(.A(n657), .B1(n651), .B2(n476), .ZN(n658));
  XNOR2_X1  g356(.A(n658), .B(n473), .ZN(n659));
  INV_X1    g357(.A(n659), .ZN(n660));
  AND3_X1   g358(.A1(625), .A2(n583), .A3(122), .ZN(n661));
  AOI221_X1 g359(.A(n661), .B1(n588), .B2(n445), .C1(n590), .C2(n660), .ZN(7470));
  OAI21_X1  g360(.A(n551), .B1(n553), .B2(n546), .ZN(n663));
  AOI211_X1 g361(.A(n651), .B(n663), .C1(n548), .C2(n547), .ZN(n664));
  XNOR2_X1  g362(.A(n664), .B(n550), .ZN(n665));
  NOR2_X1   g363(.A1(n665), .A2(n591), .ZN(n666));
  AND3_X1   g364(.A1(625), .A2(n583), .A3(128), .ZN(n667));
  AOI211_X1 g365(.A(n666), .B(n667), .C1(n588), .C2(n431), .ZN(7471));
  NOR3_X1   g366(.A1(n468), .A2(n466), .A3(n597), .ZN(n669));
  OAI21_X1  g367(.A(n553), .B1(n652), .B2(n468), .ZN(n670));
  NOR2_X1   g368(.A1(n670), .A2(n669), .ZN(n671));
  XNOR2_X1  g369(.A(n671), .B(n546), .ZN(n672));
  NOR2_X1   g370(.A1(n672), .A2(n591), .ZN(n673));
  AND3_X1   g371(.A1(625), .A2(n583), .A3(127), .ZN(n674));
  AOI211_X1 g372(.A(n673), .B(n674), .C1(n588), .C2(n438), .ZN(7472));
  OAI21_X1  g373(.A(n652), .B1(n466), .B2(n597), .ZN(n676));
  XOR2_X1   g374(.A(n676), .B(n468), .ZN(n677));
  NOR2_X1   g375(.A1(n677), .A2(n591), .ZN(n678));
  AND3_X1   g376(.A1(625), .A2(n583), .A3(126), .ZN(n679));
  AOI211_X1 g377(.A(n678), .B(n679), .C1(n588), .C2(n424), .ZN(7473));
  XOR2_X1   g378(.A(n481), .B(n479), .ZN(n681));
  XNOR2_X1  g379(.A(n485), .B(n483), .ZN(n682));
  XNOR2_X1  g380(.A(n682), .B(n681), .ZN(n683));
  XNOR2_X1  g381(.A(n494), .B(n487), .ZN(n684));
  INV_X1    g382(.A(n684), .ZN(n685));
  XOR2_X1   g383(.A(n498), .B(n491), .ZN(n686));
  MUX2_X1   g384(.S(332), .B(372), .A(369), .ZN(n687));
  XNOR2_X1  g385(.A(n687), .B(n489), .ZN(n688));
  NAND3_X1  g386(.A1(n688), .A2(n686), .A3(n685), .ZN(n689));
  OR3_X1    g387(.A1(n688), .A2(n686), .A3(n684), .ZN(n690));
  INV_X1    g388(.A(n688), .ZN(n691));
  OR3_X1    g389(.A1(n691), .A2(n686), .A3(n685), .ZN(n692));
  NAND3_X1  g390(.A1(n691), .A2(n686), .A3(n684), .ZN(n693));
  AND4_X1   g391(.A1(n692), .A2(n690), .A3(n689), .A4(n693), .ZN(n694));
  XNOR2_X1  g392(.A(n694), .B(n683), .ZN(7474));
  XOR2_X1   g393(.A(n467), .B(n465), .ZN(n696));
  XNOR2_X1  g394(.A(n475), .B(n470), .ZN(n697));
  XNOR2_X1  g395(.A(n697), .B(n696), .ZN(n698));
  XNOR2_X1  g396(.A(n472), .B(n460), .ZN(n699));
  MUX2_X1   g397(.S(335), .B(292), .A(289), .ZN(n700));
  XNOR2_X1  g398(.A(n700), .B(n455), .ZN(n701));
  INV_X1    g399(.A(n701), .ZN(n702));
  XNOR2_X1  g400(.A(n462), .B(n458), .ZN(n703));
  INV_X1    g401(.A(n703), .ZN(n704));
  NOR3_X1   g402(.A1(n704), .A2(n702), .A3(n699), .ZN(n705));
  NOR3_X1   g403(.A1(n703), .A2(n701), .A3(n699), .ZN(n706));
  INV_X1    g404(.A(n699), .ZN(n707));
  NOR3_X1   g405(.A1(n704), .A2(n701), .A3(n707), .ZN(n708));
  NOR3_X1   g406(.A1(n703), .A2(n702), .A3(n707), .ZN(n709));
  NOR4_X1   g407(.A1(n708), .A2(n706), .A3(n705), .A4(n709), .ZN(n710));
  XNOR2_X1  g408(.A(n710), .B(n698), .ZN(7476));
  INV_X1    g409(.A(n477), .ZN(n712));
  OAI21_X1  g410(.A(n559), .B1(n712), .B2(n597), .ZN(n713));
  NAND3_X1  g411(.A1(n540), .A2(n539), .A3(n459), .ZN(n714));
  OAI211_X1 g412(.A(n543), .B(n714), .C1(n537), .C2(n535), .ZN(n715));
  XNOR2_X1  g413(.A(n715), .B(n456), .ZN(n716));
  INV_X1    g414(.A(n716), .ZN(n717));
  AOI21_X1  g415(.A(n715), .B1(n464), .B2(n459), .ZN(n718));
  XNOR2_X1  g416(.A(n718), .B(n456), .ZN(n719));
  MUX2_X1   g417(.S(n713), .B(n719), .A(n717), .ZN(n720));
  INV_X1    g418(.A(n720), .ZN(n721));
  NAND4_X1  g419(.A1(n672), .A2(n665), .A3(n598), .A4(n677), .ZN(n722));
  AOI21_X1  g420(.A(n536), .B1(n540), .B2(n539), .ZN(n723));
  XNOR2_X1  g421(.A(n723), .B(n459), .ZN(n724));
  INV_X1    g422(.A(n724), .ZN(n725));
  AOI211_X1 g423(.A(n536), .B(n464), .C1(n539), .C2(n540), .ZN(n726));
  XNOR2_X1  g424(.A(n726), .B(n535), .ZN(n727));
  MUX2_X1   g425(.S(n713), .B(n727), .A(n725), .ZN(n728));
  XNOR2_X1  g426(.A(n540), .B(n539), .ZN(n729));
  NOR2_X1   g427(.A1(n460), .A2(422), .ZN(n730));
  XNOR2_X1  g428(.A(n730), .B(n539), .ZN(n731));
  INV_X1    g429(.A(n731), .ZN(n732));
  MUX2_X1   g430(.S(n713), .B(n732), .A(n729), .ZN(n733));
  INV_X1    g431(.A(n461), .ZN(n734));
  XNOR2_X1  g432(.A(n713), .B(n734), .ZN(n735));
  NAND3_X1  g433(.A1(n735), .A2(n733), .A3(n728), .ZN(n736));
  NOR4_X1   g434(.A1(n722), .A2(n721), .A3(n660), .A4(n736), .ZN(7503));
  INV_X1    g435(.A(7432), .ZN(n738));
  NAND4_X1  g436(.A1(n633), .A2(n593), .A3(n585), .A4(n640), .ZN(n739));
  AOI21_X1  g437(.A(n565), .B1(n563), .B2(n480), .ZN(n740));
  XNOR2_X1  g438(.A(n740), .B(n485), .ZN(n741));
  INV_X1    g439(.A(n741), .ZN(n742));
  AND2_X1   g440(.A1(n740), .A2(n608), .ZN(n743));
  XNOR2_X1  g441(.A(n743), .B(n562), .ZN(n744));
  MUX2_X1   g442(.S(n602), .B(n744), .A(n742), .ZN(n745));
  XNOR2_X1  g443(.A(n563), .B(n480), .ZN(n746));
  NOR2_X1   g444(.A1(n481), .A2(490), .ZN(n747));
  XNOR2_X1  g445(.A(n747), .B(n480), .ZN(n748));
  INV_X1    g446(.A(n748), .ZN(n749));
  MUX2_X1   g447(.S(n602), .B(n749), .A(n746), .ZN(n750));
  XNOR2_X1  g448(.A(n602), .B(n482), .ZN(n751));
  NAND3_X1  g449(.A1(n751), .A2(n750), .A3(n745), .ZN(n752));
  NOR4_X1   g450(.A1(n739), .A2(n629), .A3(n738), .A4(n752), .ZN(7504));
  INV_X1    g451(.A(571), .ZN(n754));
  NOR2_X1   g452(.A1(574), .A2(n754), .ZN(n755));
  INV_X1    g453(.A(n755), .ZN(n756));
  NOR2_X1   g454(.A1(574), .A2(571), .ZN(n757));
  INV_X1    g455(.A(n757), .ZN(n758));
  AND2_X1   g456(.A1(574), .A2(571), .ZN(n759));
  AND2_X1   g457(.A1(574), .A2(n754), .ZN(n760));
  AOI22_X1  g458(.A1(n759), .A2(185), .B1(182), .B2(n760), .ZN(n761));
  OAI221_X1 g459(.A(n761), .B1(n756), .B2(7365), .C1(7015), .C2(n758), .ZN(n762));
  AND2_X1   g460(.A1(n762), .A2(137), .ZN(7506));
  INV_X1    g461(.A(577), .ZN(n764));
  NOR2_X1   g462(.A1(580), .A2(n764), .ZN(n765));
  INV_X1    g463(.A(n765), .ZN(n766));
  NOR2_X1   g464(.A1(580), .A2(577), .ZN(n767));
  INV_X1    g465(.A(n767), .ZN(n768));
  NAND3_X1  g466(.A1(580), .A2(577), .A3(185), .ZN(n769));
  NAND3_X1  g467(.A1(580), .A2(n764), .A3(182), .ZN(n770));
  AND2_X1   g468(.A1(n770), .A2(n769), .ZN(n771));
  OAI221_X1 g469(.A(n771), .B1(n766), .B2(7365), .C1(7015), .C2(n768), .ZN(n772));
  AND2_X1   g470(.A1(n772), .A2(137), .ZN(7511));
  AOI22_X1  g471(.A1(n615), .A2(37), .B1(43), .B2(n616), .ZN(n774));
  OAI221_X1 g472(.A(n774), .B1(7465), .B2(n614), .C1(n613), .C2(7470), .ZN(7515));
  AOI22_X1  g473(.A1(n615), .A2(20), .B1(76), .B2(n616), .ZN(n776));
  OAI221_X1 g474(.A(n776), .B1(7466), .B2(n614), .C1(n613), .C2(7471), .ZN(7516));
  AOI22_X1  g475(.A1(n615), .A2(17), .B1(73), .B2(n616), .ZN(n778));
  OAI221_X1 g476(.A(n778), .B1(7467), .B2(n614), .C1(n613), .C2(7472), .ZN(7517));
  AOI22_X1  g477(.A1(n615), .A2(70), .B1(67), .B2(n616), .ZN(n780));
  OAI221_X1 g478(.A(n780), .B1(n614), .B2(7363), .C1(n613), .C2(7473), .ZN(7518));
  AOI22_X1  g479(.A1(n647), .A2(37), .B1(43), .B2(n648), .ZN(n782));
  OAI221_X1 g480(.A(n782), .B1(n646), .B2(7465), .C1(n645), .C2(7470), .ZN(7519));
  AOI22_X1  g481(.A1(n647), .A2(20), .B1(76), .B2(n648), .ZN(n784));
  OAI221_X1 g482(.A(n784), .B1(n646), .B2(7466), .C1(n645), .C2(7471), .ZN(7520));
  AOI22_X1  g483(.A1(n647), .A2(17), .B1(73), .B2(n648), .ZN(n786));
  OAI221_X1 g484(.A(n786), .B1(n646), .B2(7467), .C1(n645), .C2(7472), .ZN(7521));
  AOI22_X1  g485(.A1(n647), .A2(70), .B1(67), .B2(n648), .ZN(n788));
  OAI221_X1 g486(.A(n788), .B1(n646), .B2(7363), .C1(n645), .C2(7473), .ZN(7522));
  AOI22_X1  g487(.A1(n759), .A2(170), .B1(200), .B2(n760), .ZN(n790));
  OAI221_X1 g488(.A(n790), .B1(n756), .B2(7470), .C1(7465), .C2(n758), .ZN(n791));
  AND2_X1   g489(.A1(n791), .A2(137), .ZN(7600));
  AOI22_X1  g490(.A1(n759), .A2(158), .B1(188), .B2(n760), .ZN(n793));
  OAI221_X1 g491(.A(n793), .B1(n756), .B2(7473), .C1(7363), .C2(n758), .ZN(n794));
  AND2_X1   g492(.A1(n794), .A2(137), .ZN(7601));
  AOI22_X1  g493(.A1(n759), .A2(152), .B1(155), .B2(n760), .ZN(n796));
  OAI221_X1 g494(.A(n796), .B1(n756), .B2(7472), .C1(7467), .C2(n758), .ZN(n797));
  AND2_X1   g495(.A1(n797), .A2(137), .ZN(7602));
  AOI22_X1  g496(.A1(n759), .A2(146), .B1(149), .B2(n760), .ZN(n799));
  OAI221_X1 g497(.A(n799), .B1(n756), .B2(7471), .C1(7466), .C2(n758), .ZN(n800));
  AND2_X1   g498(.A1(n800), .A2(137), .ZN(7603));
  NAND3_X1  g499(.A1(580), .A2(577), .A3(170), .ZN(n802));
  NAND3_X1  g500(.A1(580), .A2(n764), .A3(200), .ZN(n803));
  AND2_X1   g501(.A1(n803), .A2(n802), .ZN(n804));
  OAI221_X1 g502(.A(n804), .B1(n766), .B2(7470), .C1(7465), .C2(n768), .ZN(n805));
  AND2_X1   g503(.A1(n805), .A2(137), .ZN(7604));
  NAND3_X1  g504(.A1(580), .A2(577), .A3(158), .ZN(n807));
  NAND3_X1  g505(.A1(580), .A2(n764), .A3(188), .ZN(n808));
  AND2_X1   g506(.A1(n808), .A2(n807), .ZN(n809));
  OAI221_X1 g507(.A(n809), .B1(n766), .B2(7473), .C1(7363), .C2(n768), .ZN(n810));
  AND2_X1   g508(.A1(n810), .A2(137), .ZN(7605));
  NAND3_X1  g509(.A1(580), .A2(577), .A3(152), .ZN(n812));
  NAND3_X1  g510(.A1(580), .A2(n764), .A3(155), .ZN(n813));
  AND2_X1   g511(.A1(n813), .A2(n812), .ZN(n814));
  OAI221_X1 g512(.A(n814), .B1(n766), .B2(7472), .C1(7467), .C2(n768), .ZN(n815));
  AND2_X1   g513(.A1(n815), .A2(137), .ZN(7606));
  NAND3_X1  g514(.A1(580), .A2(577), .A3(146), .ZN(n817));
  NAND3_X1  g515(.A1(580), .A2(n764), .A3(149), .ZN(n818));
  AND2_X1   g516(.A1(n818), .A2(n817), .ZN(n819));
  OAI221_X1 g517(.A(n819), .B1(n766), .B2(7471), .C1(7466), .C2(n768), .ZN(n820));
  AND2_X1   g518(.A1(n820), .A2(137), .ZN(7607));
  INV_X1    g519(.A(599), .ZN(n822));
  INV_X1    g520(.A(603), .ZN(n823));
  OR3_X1    g521(.A1(7432), .A2(n823), .A3(n822), .ZN(n824));
  XNOR2_X1  g522(.A(n483), .B(132), .ZN(n825));
  NOR3_X1   g523(.A1(n825), .A2(n823), .A3(599), .ZN(n826));
  INV_X1    g524(.A(123), .ZN(n827));
  NOR3_X1   g525(.A1(603), .A2(n822), .A3(n827), .ZN(n828));
  NOR3_X1   g526(.A1(n358), .A2(603), .A3(599), .ZN(n829));
  NOR3_X1   g527(.A1(n829), .A2(n828), .A3(n826), .ZN(n830));
  AOI22_X1  g528(.A1(n824), .A2(n830), .B1(631), .B2(135), .ZN(7626));
  XOR2_X1   g529(.A(n825), .B(7432), .ZN(7698));
  INV_X1    g530(.A(625), .ZN(n833));
  NOR3_X1   g531(.A1(n833), .A2(619), .A3(n827), .ZN(n834));
  AOI221_X1 g532(.A(n834), .B1(n588), .B2(n359), .C1(n590), .C2(n738), .ZN(7699));
  NOR2_X1   g533(.A1(n745), .A2(n591), .ZN(n836));
  AND3_X1   g534(.A1(625), .A2(n583), .A3(121), .ZN(n837));
  AOI211_X1 g535(.A(n836), .B(n837), .C1(n588), .C2(n354), .ZN(7700));
  NOR2_X1   g536(.A1(n750), .A2(n591), .ZN(n839));
  AND3_X1   g537(.A1(625), .A2(n583), .A3(116), .ZN(n840));
  AOI211_X1 g538(.A(n839), .B(n840), .C1(n588), .C2(n380), .ZN(7701));
  NOR2_X1   g539(.A1(n751), .A2(n591), .ZN(n842));
  AND3_X1   g540(.A1(625), .A2(n583), .A3(112), .ZN(n843));
  AOI211_X1 g541(.A(n842), .B(n843), .C1(n588), .C2(n367), .ZN(7702));
  AND4_X1   g542(.A1(556), .A2(552), .A3(386), .A4(562), .ZN(n845));
  NAND4_X1  g543(.A1(n532), .A2(559), .A3(245), .A4(n845), .ZN(n846));
  NOR4_X1   g544(.A1(7476), .A2(7474), .A3(6716), .A4(n846), .ZN(7703));
  AND3_X1   g545(.A1(625), .A2(n583), .A3(115), .ZN(n848));
  AOI221_X1 g546(.A(n848), .B1(n588), .B2(n395), .C1(n590), .C2(n721), .ZN(7704));
  NOR2_X1   g547(.A1(n728), .A2(n591), .ZN(n850));
  AND3_X1   g548(.A1(625), .A2(n583), .A3(114), .ZN(n851));
  AOI211_X1 g549(.A(n850), .B(n851), .C1(n588), .C2(n402), .ZN(7705));
  NOR2_X1   g550(.A1(n733), .A2(n591), .ZN(n853));
  AND3_X1   g551(.A1(625), .A2(n583), .A3(53), .ZN(n854));
  AOI211_X1 g552(.A(n853), .B(n854), .C1(n588), .C2(n409), .ZN(7706));
  NOR2_X1   g553(.A1(n735), .A2(n591), .ZN(n856));
  AND3_X1   g554(.A1(625), .A2(n583), .A3(113), .ZN(n857));
  AOI211_X1 g555(.A(n856), .B(n857), .C1(n588), .C2(n452), .ZN(7707));
  AOI22_X1  g556(.A1(n647), .A2(106), .B1(109), .B2(n648), .ZN(n859));
  OAI221_X1 g557(.A(n859), .B1(7699), .B2(n646), .C1(n645), .C2(7704), .ZN(7735));
  AOI22_X1  g558(.A1(n615), .A2(106), .B1(109), .B2(n616), .ZN(n861));
  OAI221_X1 g559(.A(n861), .B1(7699), .B2(n614), .C1(n613), .C2(7704), .ZN(7736));
  AOI22_X1  g560(.A1(n615), .A2(49), .B1(46), .B2(n616), .ZN(n863));
  OAI221_X1 g561(.A(n863), .B1(7700), .B2(n614), .C1(n613), .C2(7705), .ZN(7737));
  AOI22_X1  g562(.A1(n615), .A2(103), .B1(100), .B2(n616), .ZN(n865));
  OAI221_X1 g563(.A(n865), .B1(7701), .B2(n614), .C1(n613), .C2(7706), .ZN(7738));
  AOI22_X1  g564(.A1(n615), .A2(40), .B1(91), .B2(n616), .ZN(n867));
  OAI221_X1 g565(.A(n867), .B1(7702), .B2(n614), .C1(n613), .C2(7707), .ZN(7739));
  AOI22_X1  g566(.A1(n647), .A2(49), .B1(46), .B2(n648), .ZN(n869));
  OAI221_X1 g567(.A(n869), .B1(7700), .B2(n646), .C1(n645), .C2(7705), .ZN(7740));
  AOI22_X1  g568(.A1(n647), .A2(103), .B1(100), .B2(n648), .ZN(n871));
  OAI221_X1 g569(.A(n871), .B1(7701), .B2(n646), .C1(n645), .C2(7706), .ZN(7741));
  AOI22_X1  g570(.A1(n647), .A2(40), .B1(91), .B2(n648), .ZN(n873));
  OAI221_X1 g571(.A(n873), .B1(7702), .B2(n646), .C1(n645), .C2(7707), .ZN(7742));
  AOI22_X1  g572(.A1(n759), .A2(173), .B1(203), .B2(n760), .ZN(n875));
  OAI221_X1 g573(.A(n875), .B1(7702), .B2(n758), .C1(n756), .C2(7707), .ZN(n876));
  AND2_X1   g574(.A1(n876), .A2(137), .ZN(7754));
  AOI22_X1  g575(.A1(n759), .A2(167), .B1(197), .B2(n760), .ZN(n878));
  OAI221_X1 g576(.A(n878), .B1(7701), .B2(n758), .C1(n756), .C2(7706), .ZN(n879));
  AND2_X1   g577(.A1(n879), .A2(137), .ZN(7755));
  AOI22_X1  g578(.A1(n759), .A2(164), .B1(194), .B2(n760), .ZN(n881));
  OAI221_X1 g579(.A(n881), .B1(7700), .B2(n758), .C1(n756), .C2(7705), .ZN(n882));
  AND2_X1   g580(.A1(n882), .A2(137), .ZN(7756));
  AOI22_X1  g581(.A1(n759), .A2(161), .B1(191), .B2(n760), .ZN(n884));
  OAI221_X1 g582(.A(n884), .B1(7699), .B2(n758), .C1(n756), .C2(7704), .ZN(n885));
  AND2_X1   g583(.A1(n885), .A2(137), .ZN(7757));
  NAND3_X1  g584(.A1(580), .A2(577), .A3(173), .ZN(n887));
  NAND3_X1  g585(.A1(580), .A2(n764), .A3(203), .ZN(n888));
  AND2_X1   g586(.A1(n888), .A2(n887), .ZN(n889));
  OAI221_X1 g587(.A(n889), .B1(7702), .B2(n768), .C1(n766), .C2(7707), .ZN(n890));
  AND2_X1   g588(.A1(n890), .A2(137), .ZN(7758));
  NAND3_X1  g589(.A1(580), .A2(577), .A3(167), .ZN(n892));
  NAND3_X1  g590(.A1(580), .A2(n764), .A3(197), .ZN(n893));
  AND2_X1   g591(.A1(n893), .A2(n892), .ZN(n894));
  OAI221_X1 g592(.A(n894), .B1(7701), .B2(n768), .C1(n766), .C2(7706), .ZN(n895));
  AND2_X1   g593(.A1(n895), .A2(137), .ZN(7759));
  NAND3_X1  g594(.A1(580), .A2(577), .A3(164), .ZN(n897));
  NAND3_X1  g595(.A1(580), .A2(n764), .A3(194), .ZN(n898));
  AND2_X1   g596(.A1(n898), .A2(n897), .ZN(n899));
  OAI221_X1 g597(.A(n899), .B1(7700), .B2(n768), .C1(n766), .C2(7705), .ZN(n900));
  AND2_X1   g598(.A1(n900), .A2(137), .ZN(7760));
  NAND3_X1  g599(.A1(580), .A2(577), .A3(161), .ZN(n902));
  NAND3_X1  g600(.A1(580), .A2(n764), .A3(191), .ZN(n903));
  AND2_X1   g601(.A1(n903), .A2(n902), .ZN(n904));
  OAI221_X1 g602(.A(n904), .B1(7699), .B2(n768), .C1(n766), .C2(7704), .ZN(n905));
  AND2_X1   g603(.A1(n905), .A2(137), .ZN(7761));
  INV_X1    g604(.A(583), .ZN(n907));
  OR3_X1    g605(.A1(n623), .A2(n621), .A3(n569), .ZN(n908));
  XNOR2_X1  g606(.A(n908), .B(n620), .ZN(n909));
  XNOR2_X1  g607(.A(n909), .B(n638), .ZN(n910));
  XNOR2_X1  g608(.A(n910), .B(n626), .ZN(n911));
  XNOR2_X1  g609(.A(n911), .B(n489), .ZN(n912));
  XNOR2_X1  g610(.A(n912), .B(n488), .ZN(n913));
  XNOR2_X1  g611(.A(n913), .B(n492), .ZN(n914));
  XNOR2_X1  g612(.A(n914), .B(n495), .ZN(n915));
  AND2_X1   g613(.A1(n915), .A2(n499), .ZN(n916));
  OAI21_X1  g614(.A(n907), .B1(n915), .B2(n499), .ZN(n917));
  INV_X1    g615(.A(n488), .ZN(n918));
  NOR2_X1   g616(.A1(n495), .A2(n489), .ZN(n919));
  AND3_X1   g617(.A1(n919), .A2(n499), .A3(n918), .ZN(n920));
  NOR2_X1   g618(.A1(n920), .A2(n626), .ZN(n921));
  NOR2_X1   g619(.A1(n487), .A2(534), .ZN(n922));
  AOI21_X1  g620(.A(n908), .B1(n919), .B2(n918), .ZN(n923));
  XNOR2_X1  g621(.A(n923), .B(n922), .ZN(n924));
  XNOR2_X1  g622(.A(n924), .B(n921), .ZN(n925));
  XNOR2_X1  g623(.A(n925), .B(n489), .ZN(n926));
  XNOR2_X1  g624(.A(n926), .B(n488), .ZN(n927));
  XNOR2_X1  g625(.A(n927), .B(n492), .ZN(n928));
  XNOR2_X1  g626(.A(n928), .B(n495), .ZN(n929));
  XNOR2_X1  g627(.A(n929), .B(n571), .ZN(n930));
  OAI22_X1  g628(.A1(n917), .A2(n916), .B1(n907), .B2(n930), .ZN(n931));
  INV_X1    g629(.A(n480), .ZN(n932));
  XOR2_X1   g630(.A(n747), .B(n743), .ZN(n933));
  XNOR2_X1  g631(.A(n933), .B(n609), .ZN(n934));
  XOR2_X1   g632(.A(n934), .B(n482), .ZN(n935));
  XNOR2_X1  g633(.A(n935), .B(n932), .ZN(n936));
  XNOR2_X1  g634(.A(n936), .B(n561), .ZN(n937));
  XNOR2_X1  g635(.A(n937), .B(n485), .ZN(n938));
  INV_X1    g636(.A(n577), .ZN(n939));
  AND3_X1   g637(.A1(n938), .A2(n939), .A3(n907), .ZN(n940));
  AOI21_X1  g638(.A(n907), .B1(n577), .B2(n500), .ZN(n942));
  XNOR2_X1  g639(.A(n740), .B(n563), .ZN(n943));
  XOR2_X1   g640(.A(n943), .B(n605), .ZN(n944));
  XNOR2_X1  g641(.A(n944), .B(n482), .ZN(n945));
  XNOR2_X1  g642(.A(n945), .B(n932), .ZN(n946));
  XNOR2_X1  g643(.A(n946), .B(n561), .ZN(n947));
  XNOR2_X1  g644(.A(n947), .B(n562), .ZN(n948));
  AOI211_X1 g645(.A(n939), .B(n948), .C1(n503), .C2(583), .ZN(n949));
  AOI211_X1 g646(.A(n940), .B(n949), .C1(n942), .C2(n938), .ZN(n950));
  XNOR2_X1  g647(.A(n950), .B(n931), .ZN(n951));
  NAND2_X1  g648(.A1(n951), .A2(n590), .ZN(n952));
  XNOR2_X1  g649(.A(n380), .B(n367), .ZN(n953));
  XOR2_X1   g650(.A(n358), .B(n354), .ZN(n954));
  XNOR2_X1  g651(.A(n954), .B(n953), .ZN(n955));
  INV_X1    g652(.A(n352), .ZN(n956));
  AND2_X1   g653(.A1(351), .A2(242), .ZN(n957));
  AOI211_X1 g654(.A(534), .B(n957), .C1(n383), .C2(254), .ZN(n958));
  AND3_X1   g655(.A1(534), .A2(351), .A3(248), .ZN(n959));
  NOR3_X1   g656(.A1(n384), .A2(351), .A3(n350), .ZN(n960));
  NOR3_X1   g657(.A1(n960), .A2(n959), .A3(n958), .ZN(n961));
  AND2_X1   g658(.A1(341), .A2(242), .ZN(n962));
  AOI211_X1 g659(.A(523), .B(n962), .C1(n344), .C2(254), .ZN(n963));
  AND3_X1   g660(.A1(523), .A2(341), .A3(248), .ZN(n964));
  NOR3_X1   g661(.A1(n345), .A2(341), .A3(n350), .ZN(n965));
  NOR3_X1   g662(.A1(n965), .A2(n964), .A3(n963), .ZN(n966));
  XNOR2_X1  g663(.A(n966), .B(n961), .ZN(n967));
  MUX2_X1   g664(.S(514), .B(n349), .A(242), .ZN(n968));
  AND2_X1   g665(.A1(324), .A2(242), .ZN(n969));
  AOI211_X1 g666(.A(503), .B(n969), .C1(n370), .C2(254), .ZN(n970));
  AND3_X1   g667(.A1(503), .A2(324), .A3(248), .ZN(n971));
  NOR3_X1   g668(.A1(n371), .A2(324), .A3(n350), .ZN(n972));
  NOR3_X1   g669(.A1(n972), .A2(n971), .A3(n970), .ZN(n973));
  XNOR2_X1  g670(.A(n973), .B(n968), .ZN(n974));
  AND3_X1   g671(.A1(n974), .A2(n967), .A3(n956), .ZN(n975));
  NOR3_X1   g672(.A1(n974), .A2(n967), .A3(n352), .ZN(n976));
  INV_X1    g673(.A(n974), .ZN(n977));
  AND3_X1   g674(.A1(n977), .A2(n967), .A3(n352), .ZN(n978));
  NOR3_X1   g675(.A1(n977), .A2(n967), .A3(n956), .ZN(n979));
  NOR4_X1   g676(.A1(n978), .A2(n976), .A3(n975), .A4(n979), .ZN(n980));
  XNOR2_X1  g677(.A(n980), .B(n955), .ZN(n981));
  NAND2_X1  g678(.A1(n981), .A2(n588), .ZN(n982));
  OAI21_X1  g679(.A(625), .B1(619), .B2(120), .ZN(n983));
  NAND3_X1  g680(.A1(n983), .A2(n982), .A3(n952), .ZN(8075));
  INV_X1    g681(.A(566), .ZN(n985));
  OR2_X1    g682(.A1(n553), .A2(n546), .ZN(n986));
  AND3_X1   g683(.A1(n986), .A2(n653), .A3(n551), .ZN(n987));
  XNOR2_X1  g684(.A(n987), .B(n548), .ZN(n988));
  XNOR2_X1  g685(.A(n988), .B(n670), .ZN(n989));
  XNOR2_X1  g686(.A(n989), .B(n657), .ZN(n990));
  XNOR2_X1  g687(.A(n990), .B(n466), .ZN(n991));
  XNOR2_X1  g688(.A(n991), .B(n468), .ZN(n992));
  XNOR2_X1  g689(.A(n992), .B(n473), .ZN(n993));
  XNOR2_X1  g690(.A(n993), .B(n546), .ZN(n994));
  AND2_X1   g691(.A1(n994), .A2(n476), .ZN(n995));
  OAI21_X1  g692(.A(n985), .B1(n994), .B2(n476), .ZN(n996));
  NOR4_X1   g693(.A1(n546), .A2(n468), .A3(n466), .A4(n550), .ZN(n997));
  NOR2_X1   g694(.A1(n997), .A2(n657), .ZN(n998));
  NOR2_X1   g695(.A1(n670), .A2(n469), .ZN(n999));
  OR3_X1    g696(.A1(n546), .A2(n468), .A3(n466), .ZN(n1000));
  NAND4_X1  g697(.A1(n986), .A2(n653), .A3(n551), .A4(n1000), .ZN(n1001));
  NOR2_X1   g698(.A1(n465), .A2(374), .ZN(n1002));
  XNOR2_X1  g699(.A(n1002), .B(n1001), .ZN(n1003));
  XNOR2_X1  g700(.A(n1003), .B(n999), .ZN(n1004));
  XNOR2_X1  g701(.A(n1004), .B(n998), .ZN(n1005));
  XNOR2_X1  g702(.A(n1005), .B(n466), .ZN(n1006));
  XNOR2_X1  g703(.A(n1006), .B(n468), .ZN(n1007));
  XNOR2_X1  g704(.A(n1007), .B(n473), .ZN(n1008));
  XNOR2_X1  g705(.A(n1008), .B(n546), .ZN(n1009));
  XNOR2_X1  g706(.A(n1009), .B(n550), .ZN(n1010));
  OAI22_X1  g707(.A1(n996), .A2(n995), .B1(n985), .B2(n1010), .ZN(n1011));
  XOR2_X1   g708(.A(n730), .B(n726), .ZN(n1012));
  XNOR2_X1  g709(.A(n1012), .B(n718), .ZN(n1013));
  XOR2_X1   g710(.A(n1013), .B(n734), .ZN(n1014));
  XNOR2_X1  g711(.A(n1014), .B(n463), .ZN(n1015));
  XNOR2_X1  g712(.A(n1015), .B(n456), .ZN(n1016));
  XNOR2_X1  g713(.A(n1016), .B(n535), .ZN(n1017));
  NOR3_X1   g714(.A1(n1017), .A2(n559), .A3(566), .ZN(n1018));
  AOI211_X1 g715(.A(n985), .B(n1017), .C1(n559), .C2(n712), .ZN(n1019));
  INV_X1    g716(.A(n559), .ZN(n1020));
  XNOR2_X1  g717(.A(n723), .B(n540), .ZN(n1021));
  XNOR2_X1  g718(.A(n1021), .B(n715), .ZN(n1022));
  XNOR2_X1  g719(.A(n1022), .B(n461), .ZN(n1023));
  XNOR2_X1  g720(.A(n1023), .B(n463), .ZN(n1024));
  XNOR2_X1  g721(.A(n1024), .B(n456), .ZN(n1025));
  XNOR2_X1  g722(.A(n1025), .B(n535), .ZN(n1026));
  AOI211_X1 g723(.A(n1020), .B(n1026), .C1(n477), .C2(566), .ZN(n1027));
  NOR3_X1   g724(.A1(n1027), .A2(n1019), .A3(n1018), .ZN(n1028));
  XNOR2_X1  g725(.A(n1028), .B(n1011), .ZN(n1029));
  NAND2_X1  g726(.A1(n1029), .A2(n590), .ZN(n1030));
  AND2_X1   g727(.A1(242), .A2(226), .ZN(n1031));
  AOI211_X1 g728(.A(422), .B(n1031), .C1(254), .C2(n448), .ZN(n1032));
  AND3_X1   g729(.A1(422), .A2(248), .A3(226), .ZN(n1033));
  NOR3_X1   g730(.A1(n449), .A2(n350), .A3(226), .ZN(n1034));
  NOR3_X1   g731(.A1(n1034), .A2(n1033), .A3(n1032), .ZN(n1035));
  AND2_X1   g732(.A1(242), .A2(218), .ZN(n1036));
  AOI211_X1 g733(.A(468), .B(n1036), .C1(254), .C2(n405), .ZN(n1037));
  AND3_X1   g734(.A1(468), .A2(248), .A3(218), .ZN(n1038));
  NOR3_X1   g735(.A1(n406), .A2(n350), .A3(218), .ZN(n1039));
  NOR3_X1   g736(.A1(n1039), .A2(n1038), .A3(n1037), .ZN(n1040));
  XNOR2_X1  g737(.A(n1040), .B(n1035), .ZN(n1041));
  AND2_X1   g738(.A1(242), .A2(210), .ZN(n1042));
  AOI211_X1 g739(.A(457), .B(n1042), .C1(254), .C2(n398), .ZN(n1043));
  AND3_X1   g740(.A1(457), .A2(248), .A3(210), .ZN(n1044));
  NOR3_X1   g741(.A1(n399), .A2(n350), .A3(210), .ZN(n1045));
  NOR3_X1   g742(.A1(n1045), .A2(n1044), .A3(n1043), .ZN(n1046));
  XNOR2_X1  g743(.A(n1046), .B(n395), .ZN(n1047));
  XNOR2_X1  g744(.A(n1047), .B(n1041), .ZN(n1048));
  AND2_X1   g745(.A1(273), .A2(242), .ZN(n1049));
  AOI211_X1 g746(.A(411), .B(n1049), .C1(n420), .C2(254), .ZN(n1050));
  AND3_X1   g747(.A1(411), .A2(273), .A3(248), .ZN(n1051));
  NOR3_X1   g748(.A1(n421), .A2(273), .A3(n350), .ZN(n1052));
  NOR3_X1   g749(.A1(n1052), .A2(n1051), .A3(n1050), .ZN(n1053));
  AND2_X1   g750(.A1(265), .A2(242), .ZN(n1054));
  AOI211_X1 g751(.A(400), .B(n1054), .C1(n434), .C2(254), .ZN(n1055));
  AND3_X1   g752(.A1(400), .A2(265), .A3(248), .ZN(n1056));
  NOR3_X1   g753(.A1(n435), .A2(265), .A3(n350), .ZN(n1057));
  NOR3_X1   g754(.A1(n1057), .A2(n1056), .A3(n1055), .ZN(n1058));
  XNOR2_X1  g755(.A(n1058), .B(n1053), .ZN(n1059));
  AND2_X1   g756(.A1(257), .A2(242), .ZN(n1060));
  AOI211_X1 g757(.A(389), .B(n1060), .C1(n427), .C2(254), .ZN(n1061));
  AND3_X1   g758(.A1(389), .A2(257), .A3(248), .ZN(n1062));
  NOR3_X1   g759(.A1(n428), .A2(257), .A3(n350), .ZN(n1063));
  NOR3_X1   g760(.A1(n1063), .A2(n1062), .A3(n1061), .ZN(n1064));
  AND2_X1   g761(.A1(242), .A2(234), .ZN(n1065));
  AOI211_X1 g762(.A(435), .B(n1065), .C1(254), .C2(n441), .ZN(n1066));
  AND3_X1   g763(.A1(435), .A2(248), .A3(234), .ZN(n1067));
  NOR3_X1   g764(.A1(n442), .A2(n350), .A3(234), .ZN(n1068));
  NOR3_X1   g765(.A1(n1068), .A2(n1067), .A3(n1066), .ZN(n1069));
  XNOR2_X1  g766(.A(n1069), .B(n1064), .ZN(n1070));
  AND2_X1   g767(.A1(281), .A2(242), .ZN(n1071));
  AOI211_X1 g768(.A(374), .B(n1071), .C1(n413), .C2(254), .ZN(n1072));
  AND3_X1   g769(.A1(374), .A2(281), .A3(248), .ZN(n1073));
  NOR3_X1   g770(.A1(n414), .A2(281), .A3(n350), .ZN(n1074));
  NOR3_X1   g771(.A1(n1074), .A2(n1073), .A3(n1072), .ZN(n1075));
  INV_X1    g772(.A(n1075), .ZN(n1076));
  AND3_X1   g773(.A1(n1076), .A2(n1070), .A3(n1059), .ZN(n1077));
  NOR3_X1   g774(.A1(n1075), .A2(n1070), .A3(n1059), .ZN(n1078));
  INV_X1    g775(.A(n1070), .ZN(n1079));
  AND3_X1   g776(.A1(n1075), .A2(n1079), .A3(n1059), .ZN(n1080));
  NOR3_X1   g777(.A1(n1076), .A2(n1079), .A3(n1059), .ZN(n1081));
  NOR4_X1   g778(.A1(n1080), .A2(n1078), .A3(n1077), .A4(n1081), .ZN(n1082));
  XNOR2_X1  g779(.A(n1082), .B(n1048), .ZN(n1083));
  NAND2_X1  g780(.A1(n1083), .A2(n588), .ZN(n1084));
  OAI21_X1  g781(.A(625), .B1(619), .B2(118), .ZN(n1085));
  NAND3_X1  g782(.A1(n1085), .A2(n1084), .A3(n1030), .ZN(8076));
  INV_X1    g783(.A(97), .ZN(n1087));
  MUX2_X1   g784(.S(n583), .B(n1083), .A(n1029), .ZN(n1088));
  MUX2_X1   g785(.S(n833), .B(n1088), .A(n1087), .ZN(n1089));
  INV_X1    g786(.A(94), .ZN(n1090));
  MUX2_X1   g787(.S(n583), .B(n981), .A(n951), .ZN(n1091));
  MUX2_X1   g788(.S(n833), .B(n1091), .A(n1090), .ZN(n1092));
  AOI22_X1  g789(.A1(n615), .A2(64), .B1(14), .B2(n616), .ZN(n1093));
  OAI221_X1 g790(.A(n1093), .B1(n1089), .B2(n613), .C1(n614), .C2(n1092), .ZN(8123));
  AOI22_X1  g791(.A1(n647), .A2(64), .B1(14), .B2(n648), .ZN(n1095));
  OAI221_X1 g792(.A(n1095), .B1(n1089), .B2(n645), .C1(n646), .C2(n1092), .ZN(8124));
  AOI22_X1  g793(.A1(n759), .A2(179), .B1(176), .B2(n760), .ZN(n1097));
  OAI221_X1 g794(.A(n1097), .B1(n1089), .B2(n756), .C1(n758), .C2(n1092), .ZN(n1098));
  NAND2_X1  g795(.A1(n1098), .A2(137), .ZN(8127));
  AND3_X1   g796(.A1(580), .A2(577), .A3(179), .ZN(n1100));
  AND3_X1   g797(.A1(580), .A2(n764), .A3(176), .ZN(n1101));
  NOR2_X1   g798(.A1(n1101), .A2(n1100), .ZN(n1102));
  OAI221_X1 g799(.A(n1102), .B1(n1089), .B2(n766), .C1(n768), .C2(n1092), .ZN(n1103));
  NAND2_X1  g800(.A1(n1103), .A2(137), .ZN(8128));
  BUF_X1    g801(.A(141), .ZN(709));
  BUF_X1    g802(.A(293), .ZN(816));
  BUF_X1    g803(.A(592), .ZN(1066));
  INV_X1    g804(.A(545), .ZN(1142));
  INV_X1    g805(.A(545), .ZN(1143));
  BUF_X1    g806(.A(137), .ZN(2139));
  BUF_X1    g807(.A(141), .ZN(2142));
  BUF_X1    g808(.A(\1 ), .ZN(2309));
  BUF_X1    g809(.A(549), .ZN(2387));
  BUF_X1    g810(.A(299), .ZN(2527));
  INV_X1    g811(.A(549), .ZN(2584));
  BUF_X1    g812(.A(\1 ), .ZN(3357));
  BUF_X1    g813(.A(\1 ), .ZN(3358));
  BUF_X1    g814(.A(\1 ), .ZN(3359));
  BUF_X1    g815(.A(\1 ), .ZN(3360));
  BUF_X1    g816(.A(299), .ZN(3604));
  NAND3_X1  g817(.A1(n324), .A2(31), .A3(27), .ZN(4278));
endmodule


